library IEEE;
use IEEE.STD_LOGIC_1164.ALL;  
use IEEE.NUMERIC_STD.ALL;
use work.data_types.all;

entity adc is
    port (
      rst    : in std_logic;
      clk    : in std_logic;
		sndclk : out std_logic;
      data   : in std_logic;
      word   : out signed(15 downto 0)
    );
end;

architecture behavioral of adc is
  component polyphase
    Generic (
        coef_scale : integer;
        w_acc : integer;
        w_in : integer;
        w_out : integer;
        coef : array_of_integers;
        D : integer := 4
    );
    port (
      rst    : in std_logic;
      clk    : in std_logic;
      inclk : in std_logic;
      outclk : out std_logic;
      word   : in signed(w_in-1 downto 0);
      resp   : out signed(w_out-1 downto 0)
    );
  end component;



	signal interclk : std_logic := '0';
	signal input : signed(0 downto 0);
	signal inter : signed(15 downto 0);

begin
  process(clk, rst)
    variable buf : std_logic_vector(1023 downto 0);
    variable sum : unsigned(11 downto 0);
    variable data_num : unsigned(0 downto 0);
    variable last_num : unsigned(0 downto 0);
  begin
    if rst = '0' then
      buf := (others => '0');
      sum := to_unsigned(0, sum'length);
    elsif rising_edge(clk) then
	     input(0) <= data;
    end if;
  end process;
  
  filter_inst1 : polyphase
  generic map (
    coef_scale => 1,
    w_acc => 32,
    w_in => 1,
    w_out => 16,
    D => 128,
    coef => (
-29,-4,-5,-6,-5,-2,4,13,24,39,55,72,89,104,115,123,125,122,114,102,87,71,53,37,23,12,4,-2,-5,-6,-5,-4,
-3,-4,-5,-6,-4,-1,5,14,25,40,56,73,90,105,116,123,125,122,114,101,86,69,52,36,22,11,3,-2,-5,-6,-5,-4,
-3,-4,-5,-6,-4,-1,5,14,27,41,58,75,91,106,117,123,125,121,113,100,85,68,51,35,21,10,2,-3,-5,-6,-5,-4,
-3,-4,-5,-6,-4,-0,6,15,28,43,59,76,93,107,117,124,125,121,112,99,83,66,49,34,20,10,2,-3,-5,-6,-5,-4,
-3,-4,-5,-6,-4,0,7,16,29,44,61,78,94,108,118,124,125,120,111,98,82,65,48,32,19,9,1,-3,-5,-6,-5,-3,
-3,-5,-6,-5,-4,0,7,17,30,45,62,79,95,109,119,124,124,119,110,96,80,63,47,31,18,8,1,-3,-5,-6,-5,-3,
-3,-5,-6,-5,-3,1,8,18,31,47,63,80,96,110,119,124,124,119,109,95,79,62,45,30,17,7,0,-4,-5,-6,-5,-3,
-3,-5,-6,-5,-3,1,9,19,32,48,65,82,98,111,120,125,124,118,108,94,78,61,44,29,16,7,0,-4,-6,-5,-4,-3,
-4,-5,-6,-5,-3,2,10,20,34,49,66,83,99,112,121,125,124,117,107,93,76,59,43,28,15,6,-0,-4,-6,-5,-4,-3,
-4,-5,-6,-5,-3,2,10,21,35,51,68,85,100,113,121,125,123,117,106,91,75,58,41,27,14,5,-1,-4,-6,-5,-4,-3,
-4,-5,-6,-5,-2,3,11,22,36,52,69,86,101,114,122,125,123,116,105,90,73,56,40,25,14,5,-1,-4,-6,-5,-4,-3,
-4,-5,-6,-5,-2,4,12,23,37,53,71,87,102,114,122,125,123,115,104,89,72,55,39,24,13,4,-2,-5,-6,-5,-4,-29

	 )
  )
  port map (
    rst => rst,
    clk => clk,
    inclk => clk,
    outclk => interclk,
    word => input,
    resp => inter
  );
  filter_inst2 : polyphase
  generic map (
    coef_scale => 2**11,
    w_acc => 32,
    w_in => 16,
    w_out => 16,
    D => 8,
    coef => (
1,-1,1,-1,1,-1,1,0,-2,5,-9,13,-18,23,-30,41,229,11,-17,17,-16,13,-10,7,-4,2,-0,-0,1,-1,1,-1,
-0,-0,1,-1,2,-2,2,-1,-0,3,-7,12,-18,27,-40,75,219,-14,-4,10,-11,11,-9,7,-5,3,-1,0,0,-1,0,-0,
-0,-0,1,-1,2,-3,3,-3,2,0,-4,9,-16,27,-47,110,201,-33,8,2,-6,8,-8,7,-5,4,-2,1,-0,-0,0,-0,
-0,-0,0,-1,2,-3,4,-4,4,-3,0,4,-12,24,-49,144,176,-44,18,-6,-1,4,-6,6,-5,4,-3,2,-1,0,0,-0,
-0,0,0,-1,2,-3,4,-5,6,-6,4,-1,-6,18,-44,176,144,-49,24,-12,4,0,-3,4,-4,4,-3,2,-1,0,-0,-0,
-0,0,-0,-0,1,-2,4,-5,7,-8,8,-6,2,8,-33,201,110,-47,27,-16,9,-4,0,2,-3,3,-3,2,-1,1,-0,-0,
-0,0,-1,0,0,-1,3,-5,7,-9,11,-11,10,-4,-14,219,75,-40,27,-18,12,-7,3,-0,-1,2,-2,2,-1,1,-0,-0,
-1,1,-1,1,-0,-0,2,-4,7,-10,13,-16,17,-17,11,229,41,-30,23,-18,13,-9,5,-2,0,1,-1,1,-1,1,-1,1
)
  )
  port map (
    rst => rst,
    clk => clk,
    inclk => interclk,
    outclk => sndclk,
    word => inter,
    resp => word
  );


end;
