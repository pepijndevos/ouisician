-- megafunction wizard: %Shift register (RAM-based)%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTSHIFT_TAPS 

-- ============================================================
-- File Name: Shift_registers_128.vhd
-- Megafunction Name(s):
-- 			ALTSHIFT_TAPS
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 16.0.0 Build 211 04/27/2016 SJ Lite Edition
-- ************************************************************


--Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus Prime License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY Shift_registers_128 IS
	PORT
	(
		clken		: IN STD_LOGIC  := '1';
		clock		: IN STD_LOGIC ;
		shiftin		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		shiftout		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps0x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps100x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps101x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps102x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps103x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps104x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps105x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps106x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps107x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps108x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps109x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps10x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps110x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps111x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps112x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps113x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps114x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps115x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps116x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps117x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps118x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps119x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps11x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps120x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps121x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps122x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps123x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps124x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps125x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps126x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps127x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps12x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps13x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps14x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps15x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps16x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps17x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps18x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps19x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps1x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps20x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps21x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps22x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps23x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps24x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps25x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps26x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps27x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps28x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps29x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps2x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps30x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps31x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps32x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps33x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps34x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps35x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps36x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps37x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps38x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps39x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps3x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps40x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps41x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps42x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps43x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps44x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps45x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps46x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps47x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps48x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps49x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps4x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps50x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps51x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps52x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps53x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps54x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps55x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps56x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps57x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps58x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps59x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps5x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps60x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps61x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps62x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps63x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps64x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps65x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps66x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps67x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps68x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps69x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps6x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps70x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps71x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps72x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps73x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps74x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps75x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps76x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps77x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps78x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps79x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps7x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps80x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps81x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps82x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps83x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps84x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps85x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps86x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps87x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps88x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps89x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps8x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps90x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps91x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps92x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps93x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps94x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps95x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps96x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps97x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps98x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps99x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps9x		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
END Shift_registers_128;


ARCHITECTURE SYN OF shift_registers_128 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (2047 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (1615 DOWNTO 1600);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (1615 DOWNTO 1600);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (1631 DOWNTO 1616);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (1631 DOWNTO 1616);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (1647 DOWNTO 1632);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (1647 DOWNTO 1632);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (1663 DOWNTO 1648);
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (1663 DOWNTO 1648);
	SIGNAL sub_wire11	: STD_LOGIC_VECTOR (1679 DOWNTO 1664);
	SIGNAL sub_wire12	: STD_LOGIC_VECTOR (1679 DOWNTO 1664);
	SIGNAL sub_wire13	: STD_LOGIC_VECTOR (1695 DOWNTO 1680);
	SIGNAL sub_wire14	: STD_LOGIC_VECTOR (1695 DOWNTO 1680);
	SIGNAL sub_wire15	: STD_LOGIC_VECTOR (1711 DOWNTO 1696);
	SIGNAL sub_wire16	: STD_LOGIC_VECTOR (1711 DOWNTO 1696);
	SIGNAL sub_wire17	: STD_LOGIC_VECTOR (1727 DOWNTO 1712);
	SIGNAL sub_wire18	: STD_LOGIC_VECTOR (1727 DOWNTO 1712);
	SIGNAL sub_wire19	: STD_LOGIC_VECTOR (1743 DOWNTO 1728);
	SIGNAL sub_wire20	: STD_LOGIC_VECTOR (1743 DOWNTO 1728);
	SIGNAL sub_wire21	: STD_LOGIC_VECTOR (1759 DOWNTO 1744);
	SIGNAL sub_wire22	: STD_LOGIC_VECTOR (1759 DOWNTO 1744);
	SIGNAL sub_wire23	: STD_LOGIC_VECTOR (175 DOWNTO 160);
	SIGNAL sub_wire24	: STD_LOGIC_VECTOR (175 DOWNTO 160);
	SIGNAL sub_wire25	: STD_LOGIC_VECTOR (1775 DOWNTO 1760);
	SIGNAL sub_wire26	: STD_LOGIC_VECTOR (1775 DOWNTO 1760);
	SIGNAL sub_wire27	: STD_LOGIC_VECTOR (1791 DOWNTO 1776);
	SIGNAL sub_wire28	: STD_LOGIC_VECTOR (1791 DOWNTO 1776);
	SIGNAL sub_wire29	: STD_LOGIC_VECTOR (1807 DOWNTO 1792);
	SIGNAL sub_wire30	: STD_LOGIC_VECTOR (1807 DOWNTO 1792);
	SIGNAL sub_wire31	: STD_LOGIC_VECTOR (1823 DOWNTO 1808);
	SIGNAL sub_wire32	: STD_LOGIC_VECTOR (1823 DOWNTO 1808);
	SIGNAL sub_wire33	: STD_LOGIC_VECTOR (1839 DOWNTO 1824);
	SIGNAL sub_wire34	: STD_LOGIC_VECTOR (1839 DOWNTO 1824);
	SIGNAL sub_wire35	: STD_LOGIC_VECTOR (1855 DOWNTO 1840);
	SIGNAL sub_wire36	: STD_LOGIC_VECTOR (1855 DOWNTO 1840);
	SIGNAL sub_wire37	: STD_LOGIC_VECTOR (1871 DOWNTO 1856);
	SIGNAL sub_wire38	: STD_LOGIC_VECTOR (1871 DOWNTO 1856);
	SIGNAL sub_wire39	: STD_LOGIC_VECTOR (1887 DOWNTO 1872);
	SIGNAL sub_wire40	: STD_LOGIC_VECTOR (1887 DOWNTO 1872);
	SIGNAL sub_wire41	: STD_LOGIC_VECTOR (1903 DOWNTO 1888);
	SIGNAL sub_wire42	: STD_LOGIC_VECTOR (1903 DOWNTO 1888);
	SIGNAL sub_wire43	: STD_LOGIC_VECTOR (1919 DOWNTO 1904);
	SIGNAL sub_wire44	: STD_LOGIC_VECTOR (1919 DOWNTO 1904);
	SIGNAL sub_wire45	: STD_LOGIC_VECTOR (191 DOWNTO 176);
	SIGNAL sub_wire46	: STD_LOGIC_VECTOR (191 DOWNTO 176);
	SIGNAL sub_wire47	: STD_LOGIC_VECTOR (1935 DOWNTO 1920);
	SIGNAL sub_wire48	: STD_LOGIC_VECTOR (1935 DOWNTO 1920);
	SIGNAL sub_wire49	: STD_LOGIC_VECTOR (1951 DOWNTO 1936);
	SIGNAL sub_wire50	: STD_LOGIC_VECTOR (1951 DOWNTO 1936);
	SIGNAL sub_wire51	: STD_LOGIC_VECTOR (1967 DOWNTO 1952);
	SIGNAL sub_wire52	: STD_LOGIC_VECTOR (1967 DOWNTO 1952);
	SIGNAL sub_wire53	: STD_LOGIC_VECTOR (1983 DOWNTO 1968);
	SIGNAL sub_wire54	: STD_LOGIC_VECTOR (1983 DOWNTO 1968);
	SIGNAL sub_wire55	: STD_LOGIC_VECTOR (1999 DOWNTO 1984);
	SIGNAL sub_wire56	: STD_LOGIC_VECTOR (1999 DOWNTO 1984);
	SIGNAL sub_wire57	: STD_LOGIC_VECTOR (2015 DOWNTO 2000);
	SIGNAL sub_wire58	: STD_LOGIC_VECTOR (2015 DOWNTO 2000);
	SIGNAL sub_wire59	: STD_LOGIC_VECTOR (2031 DOWNTO 2016);
	SIGNAL sub_wire60	: STD_LOGIC_VECTOR (2031 DOWNTO 2016);
	SIGNAL sub_wire61	: STD_LOGIC_VECTOR (2047 DOWNTO 2032);
	SIGNAL sub_wire62	: STD_LOGIC_VECTOR (2047 DOWNTO 2032);
	SIGNAL sub_wire63	: STD_LOGIC_VECTOR (207 DOWNTO 192);
	SIGNAL sub_wire64	: STD_LOGIC_VECTOR (207 DOWNTO 192);
	SIGNAL sub_wire65	: STD_LOGIC_VECTOR (223 DOWNTO 208);
	SIGNAL sub_wire66	: STD_LOGIC_VECTOR (223 DOWNTO 208);
	SIGNAL sub_wire67	: STD_LOGIC_VECTOR (239 DOWNTO 224);
	SIGNAL sub_wire68	: STD_LOGIC_VECTOR (239 DOWNTO 224);
	SIGNAL sub_wire69	: STD_LOGIC_VECTOR (255 DOWNTO 240);
	SIGNAL sub_wire70	: STD_LOGIC_VECTOR (255 DOWNTO 240);
	SIGNAL sub_wire71	: STD_LOGIC_VECTOR (271 DOWNTO 256);
	SIGNAL sub_wire72	: STD_LOGIC_VECTOR (271 DOWNTO 256);
	SIGNAL sub_wire73	: STD_LOGIC_VECTOR (287 DOWNTO 272);
	SIGNAL sub_wire74	: STD_LOGIC_VECTOR (287 DOWNTO 272);
	SIGNAL sub_wire75	: STD_LOGIC_VECTOR (303 DOWNTO 288);
	SIGNAL sub_wire76	: STD_LOGIC_VECTOR (303 DOWNTO 288);
	SIGNAL sub_wire77	: STD_LOGIC_VECTOR (319 DOWNTO 304);
	SIGNAL sub_wire78	: STD_LOGIC_VECTOR (319 DOWNTO 304);
	SIGNAL sub_wire79	: STD_LOGIC_VECTOR (31 DOWNTO 16);
	SIGNAL sub_wire80	: STD_LOGIC_VECTOR (31 DOWNTO 16);
	SIGNAL sub_wire81	: STD_LOGIC_VECTOR (335 DOWNTO 320);
	SIGNAL sub_wire82	: STD_LOGIC_VECTOR (335 DOWNTO 320);
	SIGNAL sub_wire83	: STD_LOGIC_VECTOR (351 DOWNTO 336);
	SIGNAL sub_wire84	: STD_LOGIC_VECTOR (351 DOWNTO 336);
	SIGNAL sub_wire85	: STD_LOGIC_VECTOR (367 DOWNTO 352);
	SIGNAL sub_wire86	: STD_LOGIC_VECTOR (367 DOWNTO 352);
	SIGNAL sub_wire87	: STD_LOGIC_VECTOR (383 DOWNTO 368);
	SIGNAL sub_wire88	: STD_LOGIC_VECTOR (383 DOWNTO 368);
	SIGNAL sub_wire89	: STD_LOGIC_VECTOR (399 DOWNTO 384);
	SIGNAL sub_wire90	: STD_LOGIC_VECTOR (399 DOWNTO 384);
	SIGNAL sub_wire91	: STD_LOGIC_VECTOR (415 DOWNTO 400);
	SIGNAL sub_wire92	: STD_LOGIC_VECTOR (415 DOWNTO 400);
	SIGNAL sub_wire93	: STD_LOGIC_VECTOR (431 DOWNTO 416);
	SIGNAL sub_wire94	: STD_LOGIC_VECTOR (431 DOWNTO 416);
	SIGNAL sub_wire95	: STD_LOGIC_VECTOR (447 DOWNTO 432);
	SIGNAL sub_wire96	: STD_LOGIC_VECTOR (447 DOWNTO 432);
	SIGNAL sub_wire97	: STD_LOGIC_VECTOR (463 DOWNTO 448);
	SIGNAL sub_wire98	: STD_LOGIC_VECTOR (463 DOWNTO 448);
	SIGNAL sub_wire99	: STD_LOGIC_VECTOR (479 DOWNTO 464);
	SIGNAL sub_wire100	: STD_LOGIC_VECTOR (479 DOWNTO 464);
	SIGNAL sub_wire101	: STD_LOGIC_VECTOR (47 DOWNTO 32);
	SIGNAL sub_wire102	: STD_LOGIC_VECTOR (47 DOWNTO 32);
	SIGNAL sub_wire103	: STD_LOGIC_VECTOR (495 DOWNTO 480);
	SIGNAL sub_wire104	: STD_LOGIC_VECTOR (495 DOWNTO 480);
	SIGNAL sub_wire105	: STD_LOGIC_VECTOR (511 DOWNTO 496);
	SIGNAL sub_wire106	: STD_LOGIC_VECTOR (511 DOWNTO 496);
	SIGNAL sub_wire107	: STD_LOGIC_VECTOR (527 DOWNTO 512);
	SIGNAL sub_wire108	: STD_LOGIC_VECTOR (527 DOWNTO 512);
	SIGNAL sub_wire109	: STD_LOGIC_VECTOR (543 DOWNTO 528);
	SIGNAL sub_wire110	: STD_LOGIC_VECTOR (543 DOWNTO 528);
	SIGNAL sub_wire111	: STD_LOGIC_VECTOR (559 DOWNTO 544);
	SIGNAL sub_wire112	: STD_LOGIC_VECTOR (559 DOWNTO 544);
	SIGNAL sub_wire113	: STD_LOGIC_VECTOR (575 DOWNTO 560);
	SIGNAL sub_wire114	: STD_LOGIC_VECTOR (575 DOWNTO 560);
	SIGNAL sub_wire115	: STD_LOGIC_VECTOR (591 DOWNTO 576);
	SIGNAL sub_wire116	: STD_LOGIC_VECTOR (591 DOWNTO 576);
	SIGNAL sub_wire117	: STD_LOGIC_VECTOR (607 DOWNTO 592);
	SIGNAL sub_wire118	: STD_LOGIC_VECTOR (607 DOWNTO 592);
	SIGNAL sub_wire119	: STD_LOGIC_VECTOR (623 DOWNTO 608);
	SIGNAL sub_wire120	: STD_LOGIC_VECTOR (623 DOWNTO 608);
	SIGNAL sub_wire121	: STD_LOGIC_VECTOR (639 DOWNTO 624);
	SIGNAL sub_wire122	: STD_LOGIC_VECTOR (639 DOWNTO 624);
	SIGNAL sub_wire123	: STD_LOGIC_VECTOR (63 DOWNTO 48);
	SIGNAL sub_wire124	: STD_LOGIC_VECTOR (63 DOWNTO 48);
	SIGNAL sub_wire125	: STD_LOGIC_VECTOR (655 DOWNTO 640);
	SIGNAL sub_wire126	: STD_LOGIC_VECTOR (655 DOWNTO 640);
	SIGNAL sub_wire127	: STD_LOGIC_VECTOR (671 DOWNTO 656);
	SIGNAL sub_wire128	: STD_LOGIC_VECTOR (671 DOWNTO 656);
	SIGNAL sub_wire129	: STD_LOGIC_VECTOR (687 DOWNTO 672);
	SIGNAL sub_wire130	: STD_LOGIC_VECTOR (687 DOWNTO 672);
	SIGNAL sub_wire131	: STD_LOGIC_VECTOR (703 DOWNTO 688);
	SIGNAL sub_wire132	: STD_LOGIC_VECTOR (703 DOWNTO 688);
	SIGNAL sub_wire133	: STD_LOGIC_VECTOR (719 DOWNTO 704);
	SIGNAL sub_wire134	: STD_LOGIC_VECTOR (719 DOWNTO 704);
	SIGNAL sub_wire135	: STD_LOGIC_VECTOR (735 DOWNTO 720);
	SIGNAL sub_wire136	: STD_LOGIC_VECTOR (735 DOWNTO 720);
	SIGNAL sub_wire137	: STD_LOGIC_VECTOR (751 DOWNTO 736);
	SIGNAL sub_wire138	: STD_LOGIC_VECTOR (751 DOWNTO 736);
	SIGNAL sub_wire139	: STD_LOGIC_VECTOR (767 DOWNTO 752);
	SIGNAL sub_wire140	: STD_LOGIC_VECTOR (767 DOWNTO 752);
	SIGNAL sub_wire141	: STD_LOGIC_VECTOR (783 DOWNTO 768);
	SIGNAL sub_wire142	: STD_LOGIC_VECTOR (783 DOWNTO 768);
	SIGNAL sub_wire143	: STD_LOGIC_VECTOR (799 DOWNTO 784);
	SIGNAL sub_wire144	: STD_LOGIC_VECTOR (799 DOWNTO 784);
	SIGNAL sub_wire145	: STD_LOGIC_VECTOR (79 DOWNTO 64);
	SIGNAL sub_wire146	: STD_LOGIC_VECTOR (79 DOWNTO 64);
	SIGNAL sub_wire147	: STD_LOGIC_VECTOR (815 DOWNTO 800);
	SIGNAL sub_wire148	: STD_LOGIC_VECTOR (815 DOWNTO 800);
	SIGNAL sub_wire149	: STD_LOGIC_VECTOR (831 DOWNTO 816);
	SIGNAL sub_wire150	: STD_LOGIC_VECTOR (831 DOWNTO 816);
	SIGNAL sub_wire151	: STD_LOGIC_VECTOR (847 DOWNTO 832);
	SIGNAL sub_wire152	: STD_LOGIC_VECTOR (847 DOWNTO 832);
	SIGNAL sub_wire153	: STD_LOGIC_VECTOR (863 DOWNTO 848);
	SIGNAL sub_wire154	: STD_LOGIC_VECTOR (863 DOWNTO 848);
	SIGNAL sub_wire155	: STD_LOGIC_VECTOR (879 DOWNTO 864);
	SIGNAL sub_wire156	: STD_LOGIC_VECTOR (879 DOWNTO 864);
	SIGNAL sub_wire157	: STD_LOGIC_VECTOR (895 DOWNTO 880);
	SIGNAL sub_wire158	: STD_LOGIC_VECTOR (895 DOWNTO 880);
	SIGNAL sub_wire159	: STD_LOGIC_VECTOR (911 DOWNTO 896);
	SIGNAL sub_wire160	: STD_LOGIC_VECTOR (911 DOWNTO 896);
	SIGNAL sub_wire161	: STD_LOGIC_VECTOR (927 DOWNTO 912);
	SIGNAL sub_wire162	: STD_LOGIC_VECTOR (927 DOWNTO 912);
	SIGNAL sub_wire163	: STD_LOGIC_VECTOR (943 DOWNTO 928);
	SIGNAL sub_wire164	: STD_LOGIC_VECTOR (943 DOWNTO 928);
	SIGNAL sub_wire165	: STD_LOGIC_VECTOR (959 DOWNTO 944);
	SIGNAL sub_wire166	: STD_LOGIC_VECTOR (959 DOWNTO 944);
	SIGNAL sub_wire167	: STD_LOGIC_VECTOR (95 DOWNTO 80);
	SIGNAL sub_wire168	: STD_LOGIC_VECTOR (95 DOWNTO 80);
	SIGNAL sub_wire169	: STD_LOGIC_VECTOR (975 DOWNTO 960);
	SIGNAL sub_wire170	: STD_LOGIC_VECTOR (975 DOWNTO 960);
	SIGNAL sub_wire171	: STD_LOGIC_VECTOR (991 DOWNTO 976);
	SIGNAL sub_wire172	: STD_LOGIC_VECTOR (991 DOWNTO 976);
	SIGNAL sub_wire173	: STD_LOGIC_VECTOR (1007 DOWNTO 992);
	SIGNAL sub_wire174	: STD_LOGIC_VECTOR (1007 DOWNTO 992);
	SIGNAL sub_wire175	: STD_LOGIC_VECTOR (1023 DOWNTO 1008);
	SIGNAL sub_wire176	: STD_LOGIC_VECTOR (1023 DOWNTO 1008);
	SIGNAL sub_wire177	: STD_LOGIC_VECTOR (1039 DOWNTO 1024);
	SIGNAL sub_wire178	: STD_LOGIC_VECTOR (1039 DOWNTO 1024);
	SIGNAL sub_wire179	: STD_LOGIC_VECTOR (1055 DOWNTO 1040);
	SIGNAL sub_wire180	: STD_LOGIC_VECTOR (1055 DOWNTO 1040);
	SIGNAL sub_wire181	: STD_LOGIC_VECTOR (1071 DOWNTO 1056);
	SIGNAL sub_wire182	: STD_LOGIC_VECTOR (1071 DOWNTO 1056);
	SIGNAL sub_wire183	: STD_LOGIC_VECTOR (1087 DOWNTO 1072);
	SIGNAL sub_wire184	: STD_LOGIC_VECTOR (1087 DOWNTO 1072);
	SIGNAL sub_wire185	: STD_LOGIC_VECTOR (1103 DOWNTO 1088);
	SIGNAL sub_wire186	: STD_LOGIC_VECTOR (1103 DOWNTO 1088);
	SIGNAL sub_wire187	: STD_LOGIC_VECTOR (1119 DOWNTO 1104);
	SIGNAL sub_wire188	: STD_LOGIC_VECTOR (1119 DOWNTO 1104);
	SIGNAL sub_wire189	: STD_LOGIC_VECTOR (111 DOWNTO 96);
	SIGNAL sub_wire190	: STD_LOGIC_VECTOR (111 DOWNTO 96);
	SIGNAL sub_wire191	: STD_LOGIC_VECTOR (1135 DOWNTO 1120);
	SIGNAL sub_wire192	: STD_LOGIC_VECTOR (1135 DOWNTO 1120);
	SIGNAL sub_wire193	: STD_LOGIC_VECTOR (1151 DOWNTO 1136);
	SIGNAL sub_wire194	: STD_LOGIC_VECTOR (1151 DOWNTO 1136);
	SIGNAL sub_wire195	: STD_LOGIC_VECTOR (1167 DOWNTO 1152);
	SIGNAL sub_wire196	: STD_LOGIC_VECTOR (1167 DOWNTO 1152);
	SIGNAL sub_wire197	: STD_LOGIC_VECTOR (1183 DOWNTO 1168);
	SIGNAL sub_wire198	: STD_LOGIC_VECTOR (1183 DOWNTO 1168);
	SIGNAL sub_wire199	: STD_LOGIC_VECTOR (1199 DOWNTO 1184);
	SIGNAL sub_wire200	: STD_LOGIC_VECTOR (1199 DOWNTO 1184);
	SIGNAL sub_wire201	: STD_LOGIC_VECTOR (1215 DOWNTO 1200);
	SIGNAL sub_wire202	: STD_LOGIC_VECTOR (1215 DOWNTO 1200);
	SIGNAL sub_wire203	: STD_LOGIC_VECTOR (1231 DOWNTO 1216);
	SIGNAL sub_wire204	: STD_LOGIC_VECTOR (1231 DOWNTO 1216);
	SIGNAL sub_wire205	: STD_LOGIC_VECTOR (1247 DOWNTO 1232);
	SIGNAL sub_wire206	: STD_LOGIC_VECTOR (1247 DOWNTO 1232);
	SIGNAL sub_wire207	: STD_LOGIC_VECTOR (1263 DOWNTO 1248);
	SIGNAL sub_wire208	: STD_LOGIC_VECTOR (1263 DOWNTO 1248);
	SIGNAL sub_wire209	: STD_LOGIC_VECTOR (1279 DOWNTO 1264);
	SIGNAL sub_wire210	: STD_LOGIC_VECTOR (1279 DOWNTO 1264);
	SIGNAL sub_wire211	: STD_LOGIC_VECTOR (127 DOWNTO 112);
	SIGNAL sub_wire212	: STD_LOGIC_VECTOR (127 DOWNTO 112);
	SIGNAL sub_wire213	: STD_LOGIC_VECTOR (1295 DOWNTO 1280);
	SIGNAL sub_wire214	: STD_LOGIC_VECTOR (1295 DOWNTO 1280);
	SIGNAL sub_wire215	: STD_LOGIC_VECTOR (1311 DOWNTO 1296);
	SIGNAL sub_wire216	: STD_LOGIC_VECTOR (1311 DOWNTO 1296);
	SIGNAL sub_wire217	: STD_LOGIC_VECTOR (1327 DOWNTO 1312);
	SIGNAL sub_wire218	: STD_LOGIC_VECTOR (1327 DOWNTO 1312);
	SIGNAL sub_wire219	: STD_LOGIC_VECTOR (1343 DOWNTO 1328);
	SIGNAL sub_wire220	: STD_LOGIC_VECTOR (1343 DOWNTO 1328);
	SIGNAL sub_wire221	: STD_LOGIC_VECTOR (1359 DOWNTO 1344);
	SIGNAL sub_wire222	: STD_LOGIC_VECTOR (1359 DOWNTO 1344);
	SIGNAL sub_wire223	: STD_LOGIC_VECTOR (1375 DOWNTO 1360);
	SIGNAL sub_wire224	: STD_LOGIC_VECTOR (1375 DOWNTO 1360);
	SIGNAL sub_wire225	: STD_LOGIC_VECTOR (1391 DOWNTO 1376);
	SIGNAL sub_wire226	: STD_LOGIC_VECTOR (1391 DOWNTO 1376);
	SIGNAL sub_wire227	: STD_LOGIC_VECTOR (1407 DOWNTO 1392);
	SIGNAL sub_wire228	: STD_LOGIC_VECTOR (1407 DOWNTO 1392);
	SIGNAL sub_wire229	: STD_LOGIC_VECTOR (1423 DOWNTO 1408);
	SIGNAL sub_wire230	: STD_LOGIC_VECTOR (1423 DOWNTO 1408);
	SIGNAL sub_wire231	: STD_LOGIC_VECTOR (1439 DOWNTO 1424);
	SIGNAL sub_wire232	: STD_LOGIC_VECTOR (1439 DOWNTO 1424);
	SIGNAL sub_wire233	: STD_LOGIC_VECTOR (143 DOWNTO 128);
	SIGNAL sub_wire234	: STD_LOGIC_VECTOR (143 DOWNTO 128);
	SIGNAL sub_wire235	: STD_LOGIC_VECTOR (1455 DOWNTO 1440);
	SIGNAL sub_wire236	: STD_LOGIC_VECTOR (1455 DOWNTO 1440);
	SIGNAL sub_wire237	: STD_LOGIC_VECTOR (1471 DOWNTO 1456);
	SIGNAL sub_wire238	: STD_LOGIC_VECTOR (1471 DOWNTO 1456);
	SIGNAL sub_wire239	: STD_LOGIC_VECTOR (1487 DOWNTO 1472);
	SIGNAL sub_wire240	: STD_LOGIC_VECTOR (1487 DOWNTO 1472);
	SIGNAL sub_wire241	: STD_LOGIC_VECTOR (1503 DOWNTO 1488);
	SIGNAL sub_wire242	: STD_LOGIC_VECTOR (1503 DOWNTO 1488);
	SIGNAL sub_wire243	: STD_LOGIC_VECTOR (1519 DOWNTO 1504);
	SIGNAL sub_wire244	: STD_LOGIC_VECTOR (1519 DOWNTO 1504);
	SIGNAL sub_wire245	: STD_LOGIC_VECTOR (1535 DOWNTO 1520);
	SIGNAL sub_wire246	: STD_LOGIC_VECTOR (1535 DOWNTO 1520);
	SIGNAL sub_wire247	: STD_LOGIC_VECTOR (1551 DOWNTO 1536);
	SIGNAL sub_wire248	: STD_LOGIC_VECTOR (1551 DOWNTO 1536);
	SIGNAL sub_wire249	: STD_LOGIC_VECTOR (1567 DOWNTO 1552);
	SIGNAL sub_wire250	: STD_LOGIC_VECTOR (1567 DOWNTO 1552);
	SIGNAL sub_wire251	: STD_LOGIC_VECTOR (1583 DOWNTO 1568);
	SIGNAL sub_wire252	: STD_LOGIC_VECTOR (1583 DOWNTO 1568);
	SIGNAL sub_wire253	: STD_LOGIC_VECTOR (1599 DOWNTO 1584);
	SIGNAL sub_wire254	: STD_LOGIC_VECTOR (1599 DOWNTO 1584);
	SIGNAL sub_wire255	: STD_LOGIC_VECTOR (159 DOWNTO 144);



	COMPONENT altshift_taps
	GENERIC (
		intended_device_family		: STRING;
		lpm_hint		: STRING;
		lpm_type		: STRING;
		number_of_taps		: NATURAL;
		tap_distance		: NATURAL;
		width		: NATURAL
	);
	PORT (
			clken	: IN STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			shiftin	: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			shiftout	: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			taps	: OUT STD_LOGIC_VECTOR (2047 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	shiftout    <= sub_wire0(15 DOWNTO 0);
	sub_wire255    <= sub_wire1(159 DOWNTO 144);
	sub_wire254    <= sub_wire1(1599 DOWNTO 1584);
	sub_wire253    <= sub_wire254(1599 DOWNTO 1584);
	sub_wire252    <= sub_wire1(1583 DOWNTO 1568);
	sub_wire251    <= sub_wire252(1583 DOWNTO 1568);
	sub_wire250    <= sub_wire1(1567 DOWNTO 1552);
	sub_wire249    <= sub_wire250(1567 DOWNTO 1552);
	sub_wire248    <= sub_wire1(1551 DOWNTO 1536);
	sub_wire247    <= sub_wire248(1551 DOWNTO 1536);
	sub_wire246    <= sub_wire1(1535 DOWNTO 1520);
	sub_wire245    <= sub_wire246(1535 DOWNTO 1520);
	sub_wire244    <= sub_wire1(1519 DOWNTO 1504);
	sub_wire243    <= sub_wire244(1519 DOWNTO 1504);
	sub_wire242    <= sub_wire1(1503 DOWNTO 1488);
	sub_wire241    <= sub_wire242(1503 DOWNTO 1488);
	sub_wire240    <= sub_wire1(1487 DOWNTO 1472);
	sub_wire239    <= sub_wire240(1487 DOWNTO 1472);
	sub_wire238    <= sub_wire1(1471 DOWNTO 1456);
	sub_wire237    <= sub_wire238(1471 DOWNTO 1456);
	sub_wire236    <= sub_wire1(1455 DOWNTO 1440);
	sub_wire235    <= sub_wire236(1455 DOWNTO 1440);
	sub_wire234    <= sub_wire1(143 DOWNTO 128);
	sub_wire233    <= sub_wire234(143 DOWNTO 128);
	sub_wire232    <= sub_wire1(1439 DOWNTO 1424);
	sub_wire231    <= sub_wire232(1439 DOWNTO 1424);
	sub_wire230    <= sub_wire1(1423 DOWNTO 1408);
	sub_wire229    <= sub_wire230(1423 DOWNTO 1408);
	sub_wire228    <= sub_wire1(1407 DOWNTO 1392);
	sub_wire227    <= sub_wire228(1407 DOWNTO 1392);
	sub_wire226    <= sub_wire1(1391 DOWNTO 1376);
	sub_wire225    <= sub_wire226(1391 DOWNTO 1376);
	sub_wire224    <= sub_wire1(1375 DOWNTO 1360);
	sub_wire223    <= sub_wire224(1375 DOWNTO 1360);
	sub_wire222    <= sub_wire1(1359 DOWNTO 1344);
	sub_wire221    <= sub_wire222(1359 DOWNTO 1344);
	sub_wire220    <= sub_wire1(1343 DOWNTO 1328);
	sub_wire219    <= sub_wire220(1343 DOWNTO 1328);
	sub_wire218    <= sub_wire1(1327 DOWNTO 1312);
	sub_wire217    <= sub_wire218(1327 DOWNTO 1312);
	sub_wire216    <= sub_wire1(1311 DOWNTO 1296);
	sub_wire215    <= sub_wire216(1311 DOWNTO 1296);
	sub_wire214    <= sub_wire1(1295 DOWNTO 1280);
	sub_wire213    <= sub_wire214(1295 DOWNTO 1280);
	sub_wire212    <= sub_wire1(127 DOWNTO 112);
	sub_wire211    <= sub_wire212(127 DOWNTO 112);
	sub_wire210    <= sub_wire1(1279 DOWNTO 1264);
	sub_wire209    <= sub_wire210(1279 DOWNTO 1264);
	sub_wire208    <= sub_wire1(1263 DOWNTO 1248);
	sub_wire207    <= sub_wire208(1263 DOWNTO 1248);
	sub_wire206    <= sub_wire1(1247 DOWNTO 1232);
	sub_wire205    <= sub_wire206(1247 DOWNTO 1232);
	sub_wire204    <= sub_wire1(1231 DOWNTO 1216);
	sub_wire203    <= sub_wire204(1231 DOWNTO 1216);
	sub_wire202    <= sub_wire1(1215 DOWNTO 1200);
	sub_wire201    <= sub_wire202(1215 DOWNTO 1200);
	sub_wire200    <= sub_wire1(1199 DOWNTO 1184);
	sub_wire199    <= sub_wire200(1199 DOWNTO 1184);
	sub_wire198    <= sub_wire1(1183 DOWNTO 1168);
	sub_wire197    <= sub_wire198(1183 DOWNTO 1168);
	sub_wire196    <= sub_wire1(1167 DOWNTO 1152);
	sub_wire195    <= sub_wire196(1167 DOWNTO 1152);
	sub_wire194    <= sub_wire1(1151 DOWNTO 1136);
	sub_wire193    <= sub_wire194(1151 DOWNTO 1136);
	sub_wire192    <= sub_wire1(1135 DOWNTO 1120);
	sub_wire191    <= sub_wire192(1135 DOWNTO 1120);
	sub_wire190    <= sub_wire1(111 DOWNTO 96);
	sub_wire189    <= sub_wire190(111 DOWNTO 96);
	sub_wire188    <= sub_wire1(1119 DOWNTO 1104);
	sub_wire187    <= sub_wire188(1119 DOWNTO 1104);
	sub_wire186    <= sub_wire1(1103 DOWNTO 1088);
	sub_wire185    <= sub_wire186(1103 DOWNTO 1088);
	sub_wire184    <= sub_wire1(1087 DOWNTO 1072);
	sub_wire183    <= sub_wire184(1087 DOWNTO 1072);
	sub_wire182    <= sub_wire1(1071 DOWNTO 1056);
	sub_wire181    <= sub_wire182(1071 DOWNTO 1056);
	sub_wire180    <= sub_wire1(1055 DOWNTO 1040);
	sub_wire179    <= sub_wire180(1055 DOWNTO 1040);
	sub_wire178    <= sub_wire1(1039 DOWNTO 1024);
	sub_wire177    <= sub_wire178(1039 DOWNTO 1024);
	sub_wire176    <= sub_wire1(1023 DOWNTO 1008);
	sub_wire175    <= sub_wire176(1023 DOWNTO 1008);
	sub_wire174    <= sub_wire1(1007 DOWNTO 992);
	sub_wire173    <= sub_wire174(1007 DOWNTO 992);
	sub_wire172    <= sub_wire1(991 DOWNTO 976);
	sub_wire171    <= sub_wire172(991 DOWNTO 976);
	sub_wire170    <= sub_wire1(975 DOWNTO 960);
	sub_wire169    <= sub_wire170(975 DOWNTO 960);
	sub_wire168    <= sub_wire1(95 DOWNTO 80);
	sub_wire167    <= sub_wire168(95 DOWNTO 80);
	sub_wire166    <= sub_wire1(959 DOWNTO 944);
	sub_wire165    <= sub_wire166(959 DOWNTO 944);
	sub_wire164    <= sub_wire1(943 DOWNTO 928);
	sub_wire163    <= sub_wire164(943 DOWNTO 928);
	sub_wire162    <= sub_wire1(927 DOWNTO 912);
	sub_wire161    <= sub_wire162(927 DOWNTO 912);
	sub_wire160    <= sub_wire1(911 DOWNTO 896);
	sub_wire159    <= sub_wire160(911 DOWNTO 896);
	sub_wire158    <= sub_wire1(895 DOWNTO 880);
	sub_wire157    <= sub_wire158(895 DOWNTO 880);
	sub_wire156    <= sub_wire1(879 DOWNTO 864);
	sub_wire155    <= sub_wire156(879 DOWNTO 864);
	sub_wire154    <= sub_wire1(863 DOWNTO 848);
	sub_wire153    <= sub_wire154(863 DOWNTO 848);
	sub_wire152    <= sub_wire1(847 DOWNTO 832);
	sub_wire151    <= sub_wire152(847 DOWNTO 832);
	sub_wire150    <= sub_wire1(831 DOWNTO 816);
	sub_wire149    <= sub_wire150(831 DOWNTO 816);
	sub_wire148    <= sub_wire1(815 DOWNTO 800);
	sub_wire147    <= sub_wire148(815 DOWNTO 800);
	sub_wire146    <= sub_wire1(79 DOWNTO 64);
	sub_wire145    <= sub_wire146(79 DOWNTO 64);
	sub_wire144    <= sub_wire1(799 DOWNTO 784);
	sub_wire143    <= sub_wire144(799 DOWNTO 784);
	sub_wire142    <= sub_wire1(783 DOWNTO 768);
	sub_wire141    <= sub_wire142(783 DOWNTO 768);
	sub_wire140    <= sub_wire1(767 DOWNTO 752);
	sub_wire139    <= sub_wire140(767 DOWNTO 752);
	sub_wire138    <= sub_wire1(751 DOWNTO 736);
	sub_wire137    <= sub_wire138(751 DOWNTO 736);
	sub_wire136    <= sub_wire1(735 DOWNTO 720);
	sub_wire135    <= sub_wire136(735 DOWNTO 720);
	sub_wire134    <= sub_wire1(719 DOWNTO 704);
	sub_wire133    <= sub_wire134(719 DOWNTO 704);
	sub_wire132    <= sub_wire1(703 DOWNTO 688);
	sub_wire131    <= sub_wire132(703 DOWNTO 688);
	sub_wire130    <= sub_wire1(687 DOWNTO 672);
	sub_wire129    <= sub_wire130(687 DOWNTO 672);
	sub_wire128    <= sub_wire1(671 DOWNTO 656);
	sub_wire127    <= sub_wire128(671 DOWNTO 656);
	sub_wire126    <= sub_wire1(655 DOWNTO 640);
	sub_wire125    <= sub_wire126(655 DOWNTO 640);
	sub_wire124    <= sub_wire1(63 DOWNTO 48);
	sub_wire123    <= sub_wire124(63 DOWNTO 48);
	sub_wire122    <= sub_wire1(639 DOWNTO 624);
	sub_wire121    <= sub_wire122(639 DOWNTO 624);
	sub_wire120    <= sub_wire1(623 DOWNTO 608);
	sub_wire119    <= sub_wire120(623 DOWNTO 608);
	sub_wire118    <= sub_wire1(607 DOWNTO 592);
	sub_wire117    <= sub_wire118(607 DOWNTO 592);
	sub_wire116    <= sub_wire1(591 DOWNTO 576);
	sub_wire115    <= sub_wire116(591 DOWNTO 576);
	sub_wire114    <= sub_wire1(575 DOWNTO 560);
	sub_wire113    <= sub_wire114(575 DOWNTO 560);
	sub_wire112    <= sub_wire1(559 DOWNTO 544);
	sub_wire111    <= sub_wire112(559 DOWNTO 544);
	sub_wire110    <= sub_wire1(543 DOWNTO 528);
	sub_wire109    <= sub_wire110(543 DOWNTO 528);
	sub_wire108    <= sub_wire1(527 DOWNTO 512);
	sub_wire107    <= sub_wire108(527 DOWNTO 512);
	sub_wire106    <= sub_wire1(511 DOWNTO 496);
	sub_wire105    <= sub_wire106(511 DOWNTO 496);
	sub_wire104    <= sub_wire1(495 DOWNTO 480);
	sub_wire103    <= sub_wire104(495 DOWNTO 480);
	sub_wire102    <= sub_wire1(47 DOWNTO 32);
	sub_wire101    <= sub_wire102(47 DOWNTO 32);
	sub_wire100    <= sub_wire1(479 DOWNTO 464);
	sub_wire99    <= sub_wire100(479 DOWNTO 464);
	sub_wire98    <= sub_wire1(463 DOWNTO 448);
	sub_wire97    <= sub_wire98(463 DOWNTO 448);
	sub_wire96    <= sub_wire1(447 DOWNTO 432);
	sub_wire95    <= sub_wire96(447 DOWNTO 432);
	sub_wire94    <= sub_wire1(431 DOWNTO 416);
	sub_wire93    <= sub_wire94(431 DOWNTO 416);
	sub_wire92    <= sub_wire1(415 DOWNTO 400);
	sub_wire91    <= sub_wire92(415 DOWNTO 400);
	sub_wire90    <= sub_wire1(399 DOWNTO 384);
	sub_wire89    <= sub_wire90(399 DOWNTO 384);
	sub_wire88    <= sub_wire1(383 DOWNTO 368);
	sub_wire87    <= sub_wire88(383 DOWNTO 368);
	sub_wire86    <= sub_wire1(367 DOWNTO 352);
	sub_wire85    <= sub_wire86(367 DOWNTO 352);
	sub_wire84    <= sub_wire1(351 DOWNTO 336);
	sub_wire83    <= sub_wire84(351 DOWNTO 336);
	sub_wire82    <= sub_wire1(335 DOWNTO 320);
	sub_wire81    <= sub_wire82(335 DOWNTO 320);
	sub_wire80    <= sub_wire1(31 DOWNTO 16);
	sub_wire79    <= sub_wire80(31 DOWNTO 16);
	sub_wire78    <= sub_wire1(319 DOWNTO 304);
	sub_wire77    <= sub_wire78(319 DOWNTO 304);
	sub_wire76    <= sub_wire1(303 DOWNTO 288);
	sub_wire75    <= sub_wire76(303 DOWNTO 288);
	sub_wire74    <= sub_wire1(287 DOWNTO 272);
	sub_wire73    <= sub_wire74(287 DOWNTO 272);
	sub_wire72    <= sub_wire1(271 DOWNTO 256);
	sub_wire71    <= sub_wire72(271 DOWNTO 256);
	sub_wire70    <= sub_wire1(255 DOWNTO 240);
	sub_wire69    <= sub_wire70(255 DOWNTO 240);
	sub_wire68    <= sub_wire1(239 DOWNTO 224);
	sub_wire67    <= sub_wire68(239 DOWNTO 224);
	sub_wire66    <= sub_wire1(223 DOWNTO 208);
	sub_wire65    <= sub_wire66(223 DOWNTO 208);
	sub_wire64    <= sub_wire1(207 DOWNTO 192);
	sub_wire63    <= sub_wire64(207 DOWNTO 192);
	sub_wire62    <= sub_wire1(2047 DOWNTO 2032);
	sub_wire61    <= sub_wire62(2047 DOWNTO 2032);
	sub_wire60    <= sub_wire1(2031 DOWNTO 2016);
	sub_wire59    <= sub_wire60(2031 DOWNTO 2016);
	sub_wire58    <= sub_wire1(2015 DOWNTO 2000);
	sub_wire57    <= sub_wire58(2015 DOWNTO 2000);
	sub_wire56    <= sub_wire1(1999 DOWNTO 1984);
	sub_wire55    <= sub_wire56(1999 DOWNTO 1984);
	sub_wire54    <= sub_wire1(1983 DOWNTO 1968);
	sub_wire53    <= sub_wire54(1983 DOWNTO 1968);
	sub_wire52    <= sub_wire1(1967 DOWNTO 1952);
	sub_wire51    <= sub_wire52(1967 DOWNTO 1952);
	sub_wire50    <= sub_wire1(1951 DOWNTO 1936);
	sub_wire49    <= sub_wire50(1951 DOWNTO 1936);
	sub_wire48    <= sub_wire1(1935 DOWNTO 1920);
	sub_wire47    <= sub_wire48(1935 DOWNTO 1920);
	sub_wire46    <= sub_wire1(191 DOWNTO 176);
	sub_wire45    <= sub_wire46(191 DOWNTO 176);
	sub_wire44    <= sub_wire1(1919 DOWNTO 1904);
	sub_wire43    <= sub_wire44(1919 DOWNTO 1904);
	sub_wire42    <= sub_wire1(1903 DOWNTO 1888);
	sub_wire41    <= sub_wire42(1903 DOWNTO 1888);
	sub_wire40    <= sub_wire1(1887 DOWNTO 1872);
	sub_wire39    <= sub_wire40(1887 DOWNTO 1872);
	sub_wire38    <= sub_wire1(1871 DOWNTO 1856);
	sub_wire37    <= sub_wire38(1871 DOWNTO 1856);
	sub_wire36    <= sub_wire1(1855 DOWNTO 1840);
	sub_wire35    <= sub_wire36(1855 DOWNTO 1840);
	sub_wire34    <= sub_wire1(1839 DOWNTO 1824);
	sub_wire33    <= sub_wire34(1839 DOWNTO 1824);
	sub_wire32    <= sub_wire1(1823 DOWNTO 1808);
	sub_wire31    <= sub_wire32(1823 DOWNTO 1808);
	sub_wire30    <= sub_wire1(1807 DOWNTO 1792);
	sub_wire29    <= sub_wire30(1807 DOWNTO 1792);
	sub_wire28    <= sub_wire1(1791 DOWNTO 1776);
	sub_wire27    <= sub_wire28(1791 DOWNTO 1776);
	sub_wire26    <= sub_wire1(1775 DOWNTO 1760);
	sub_wire25    <= sub_wire26(1775 DOWNTO 1760);
	sub_wire24    <= sub_wire1(175 DOWNTO 160);
	sub_wire23    <= sub_wire24(175 DOWNTO 160);
	sub_wire22    <= sub_wire1(1759 DOWNTO 1744);
	sub_wire21    <= sub_wire22(1759 DOWNTO 1744);
	sub_wire20    <= sub_wire1(1743 DOWNTO 1728);
	sub_wire19    <= sub_wire20(1743 DOWNTO 1728);
	sub_wire18    <= sub_wire1(1727 DOWNTO 1712);
	sub_wire17    <= sub_wire18(1727 DOWNTO 1712);
	sub_wire16    <= sub_wire1(1711 DOWNTO 1696);
	sub_wire15    <= sub_wire16(1711 DOWNTO 1696);
	sub_wire14    <= sub_wire1(1695 DOWNTO 1680);
	sub_wire13    <= sub_wire14(1695 DOWNTO 1680);
	sub_wire12    <= sub_wire1(1679 DOWNTO 1664);
	sub_wire11    <= sub_wire12(1679 DOWNTO 1664);
	sub_wire10    <= sub_wire1(1663 DOWNTO 1648);
	sub_wire9    <= sub_wire10(1663 DOWNTO 1648);
	sub_wire8    <= sub_wire1(1647 DOWNTO 1632);
	sub_wire7    <= sub_wire8(1647 DOWNTO 1632);
	sub_wire6    <= sub_wire1(1631 DOWNTO 1616);
	sub_wire5    <= sub_wire6(1631 DOWNTO 1616);
	sub_wire4    <= sub_wire1(1615 DOWNTO 1600);
	sub_wire3    <= sub_wire4(1615 DOWNTO 1600);
	sub_wire2    <= sub_wire1(15 DOWNTO 0);
	taps0x    <= sub_wire2(15 DOWNTO 0);
	taps100x    <= sub_wire3(1615 DOWNTO 1600);
	taps101x    <= sub_wire5(1631 DOWNTO 1616);
	taps102x    <= sub_wire7(1647 DOWNTO 1632);
	taps103x    <= sub_wire9(1663 DOWNTO 1648);
	taps104x    <= sub_wire11(1679 DOWNTO 1664);
	taps105x    <= sub_wire13(1695 DOWNTO 1680);
	taps106x    <= sub_wire15(1711 DOWNTO 1696);
	taps107x    <= sub_wire17(1727 DOWNTO 1712);
	taps108x    <= sub_wire19(1743 DOWNTO 1728);
	taps109x    <= sub_wire21(1759 DOWNTO 1744);
	taps10x    <= sub_wire23(175 DOWNTO 160);
	taps110x    <= sub_wire25(1775 DOWNTO 1760);
	taps111x    <= sub_wire27(1791 DOWNTO 1776);
	taps112x    <= sub_wire29(1807 DOWNTO 1792);
	taps113x    <= sub_wire31(1823 DOWNTO 1808);
	taps114x    <= sub_wire33(1839 DOWNTO 1824);
	taps115x    <= sub_wire35(1855 DOWNTO 1840);
	taps116x    <= sub_wire37(1871 DOWNTO 1856);
	taps117x    <= sub_wire39(1887 DOWNTO 1872);
	taps118x    <= sub_wire41(1903 DOWNTO 1888);
	taps119x    <= sub_wire43(1919 DOWNTO 1904);
	taps11x    <= sub_wire45(191 DOWNTO 176);
	taps120x    <= sub_wire47(1935 DOWNTO 1920);
	taps121x    <= sub_wire49(1951 DOWNTO 1936);
	taps122x    <= sub_wire51(1967 DOWNTO 1952);
	taps123x    <= sub_wire53(1983 DOWNTO 1968);
	taps124x    <= sub_wire55(1999 DOWNTO 1984);
	taps125x    <= sub_wire57(2015 DOWNTO 2000);
	taps126x    <= sub_wire59(2031 DOWNTO 2016);
	taps127x    <= sub_wire61(2047 DOWNTO 2032);
	taps12x    <= sub_wire63(207 DOWNTO 192);
	taps13x    <= sub_wire65(223 DOWNTO 208);
	taps14x    <= sub_wire67(239 DOWNTO 224);
	taps15x    <= sub_wire69(255 DOWNTO 240);
	taps16x    <= sub_wire71(271 DOWNTO 256);
	taps17x    <= sub_wire73(287 DOWNTO 272);
	taps18x    <= sub_wire75(303 DOWNTO 288);
	taps19x    <= sub_wire77(319 DOWNTO 304);
	taps1x    <= sub_wire79(31 DOWNTO 16);
	taps20x    <= sub_wire81(335 DOWNTO 320);
	taps21x    <= sub_wire83(351 DOWNTO 336);
	taps22x    <= sub_wire85(367 DOWNTO 352);
	taps23x    <= sub_wire87(383 DOWNTO 368);
	taps24x    <= sub_wire89(399 DOWNTO 384);
	taps25x    <= sub_wire91(415 DOWNTO 400);
	taps26x    <= sub_wire93(431 DOWNTO 416);
	taps27x    <= sub_wire95(447 DOWNTO 432);
	taps28x    <= sub_wire97(463 DOWNTO 448);
	taps29x    <= sub_wire99(479 DOWNTO 464);
	taps2x    <= sub_wire101(47 DOWNTO 32);
	taps30x    <= sub_wire103(495 DOWNTO 480);
	taps31x    <= sub_wire105(511 DOWNTO 496);
	taps32x    <= sub_wire107(527 DOWNTO 512);
	taps33x    <= sub_wire109(543 DOWNTO 528);
	taps34x    <= sub_wire111(559 DOWNTO 544);
	taps35x    <= sub_wire113(575 DOWNTO 560);
	taps36x    <= sub_wire115(591 DOWNTO 576);
	taps37x    <= sub_wire117(607 DOWNTO 592);
	taps38x    <= sub_wire119(623 DOWNTO 608);
	taps39x    <= sub_wire121(639 DOWNTO 624);
	taps3x    <= sub_wire123(63 DOWNTO 48);
	taps40x    <= sub_wire125(655 DOWNTO 640);
	taps41x    <= sub_wire127(671 DOWNTO 656);
	taps42x    <= sub_wire129(687 DOWNTO 672);
	taps43x    <= sub_wire131(703 DOWNTO 688);
	taps44x    <= sub_wire133(719 DOWNTO 704);
	taps45x    <= sub_wire135(735 DOWNTO 720);
	taps46x    <= sub_wire137(751 DOWNTO 736);
	taps47x    <= sub_wire139(767 DOWNTO 752);
	taps48x    <= sub_wire141(783 DOWNTO 768);
	taps49x    <= sub_wire143(799 DOWNTO 784);
	taps4x    <= sub_wire145(79 DOWNTO 64);
	taps50x    <= sub_wire147(815 DOWNTO 800);
	taps51x    <= sub_wire149(831 DOWNTO 816);
	taps52x    <= sub_wire151(847 DOWNTO 832);
	taps53x    <= sub_wire153(863 DOWNTO 848);
	taps54x    <= sub_wire155(879 DOWNTO 864);
	taps55x    <= sub_wire157(895 DOWNTO 880);
	taps56x    <= sub_wire159(911 DOWNTO 896);
	taps57x    <= sub_wire161(927 DOWNTO 912);
	taps58x    <= sub_wire163(943 DOWNTO 928);
	taps59x    <= sub_wire165(959 DOWNTO 944);
	taps5x    <= sub_wire167(95 DOWNTO 80);
	taps60x    <= sub_wire169(975 DOWNTO 960);
	taps61x    <= sub_wire171(991 DOWNTO 976);
	taps62x    <= sub_wire173(1007 DOWNTO 992);
	taps63x    <= sub_wire175(1023 DOWNTO 1008);
	taps64x    <= sub_wire177(1039 DOWNTO 1024);
	taps65x    <= sub_wire179(1055 DOWNTO 1040);
	taps66x    <= sub_wire181(1071 DOWNTO 1056);
	taps67x    <= sub_wire183(1087 DOWNTO 1072);
	taps68x    <= sub_wire185(1103 DOWNTO 1088);
	taps69x    <= sub_wire187(1119 DOWNTO 1104);
	taps6x    <= sub_wire189(111 DOWNTO 96);
	taps70x    <= sub_wire191(1135 DOWNTO 1120);
	taps71x    <= sub_wire193(1151 DOWNTO 1136);
	taps72x    <= sub_wire195(1167 DOWNTO 1152);
	taps73x    <= sub_wire197(1183 DOWNTO 1168);
	taps74x    <= sub_wire199(1199 DOWNTO 1184);
	taps75x    <= sub_wire201(1215 DOWNTO 1200);
	taps76x    <= sub_wire203(1231 DOWNTO 1216);
	taps77x    <= sub_wire205(1247 DOWNTO 1232);
	taps78x    <= sub_wire207(1263 DOWNTO 1248);
	taps79x    <= sub_wire209(1279 DOWNTO 1264);
	taps7x    <= sub_wire211(127 DOWNTO 112);
	taps80x    <= sub_wire213(1295 DOWNTO 1280);
	taps81x    <= sub_wire215(1311 DOWNTO 1296);
	taps82x    <= sub_wire217(1327 DOWNTO 1312);
	taps83x    <= sub_wire219(1343 DOWNTO 1328);
	taps84x    <= sub_wire221(1359 DOWNTO 1344);
	taps85x    <= sub_wire223(1375 DOWNTO 1360);
	taps86x    <= sub_wire225(1391 DOWNTO 1376);
	taps87x    <= sub_wire227(1407 DOWNTO 1392);
	taps88x    <= sub_wire229(1423 DOWNTO 1408);
	taps89x    <= sub_wire231(1439 DOWNTO 1424);
	taps8x    <= sub_wire233(143 DOWNTO 128);
	taps90x    <= sub_wire235(1455 DOWNTO 1440);
	taps91x    <= sub_wire237(1471 DOWNTO 1456);
	taps92x    <= sub_wire239(1487 DOWNTO 1472);
	taps93x    <= sub_wire241(1503 DOWNTO 1488);
	taps94x    <= sub_wire243(1519 DOWNTO 1504);
	taps95x    <= sub_wire245(1535 DOWNTO 1520);
	taps96x    <= sub_wire247(1551 DOWNTO 1536);
	taps97x    <= sub_wire249(1567 DOWNTO 1552);
	taps98x    <= sub_wire251(1583 DOWNTO 1568);
	taps99x    <= sub_wire253(1599 DOWNTO 1584);
	taps9x    <= sub_wire255(159 DOWNTO 144);

	ALTSHIFT_TAPS_component : ALTSHIFT_TAPS
	GENERIC MAP (
		intended_device_family => "Cyclone V",
		lpm_hint => "RAM_BLOCK_TYPE=M10K",
		lpm_type => "altshift_taps",
		number_of_taps => 128,
		tap_distance => 16,
		width => 16
	)
	PORT MAP (
		clken => clken,
		clock => clock,
		shiftin => shiftin,
		shiftout => sub_wire0,
		taps => sub_wire1
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ACLR NUMERIC "0"
-- Retrieval info: PRIVATE: CLKEN NUMERIC "1"
-- Retrieval info: PRIVATE: GROUP_TAPS NUMERIC "1"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: PRIVATE: NUMBER_OF_TAPS NUMERIC "128"
-- Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: TAP_DISTANCE NUMERIC "16"
-- Retrieval info: PRIVATE: WIDTH NUMERIC "16"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: LPM_HINT STRING "RAM_BLOCK_TYPE=M10K"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altshift_taps"
-- Retrieval info: CONSTANT: NUMBER_OF_TAPS NUMERIC "128"
-- Retrieval info: CONSTANT: TAP_DISTANCE NUMERIC "16"
-- Retrieval info: CONSTANT: WIDTH NUMERIC "16"
-- Retrieval info: USED_PORT: clken 0 0 0 0 INPUT VCC "clken"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: shiftin 0 0 16 0 INPUT NODEFVAL "shiftin[15..0]"
-- Retrieval info: USED_PORT: shiftout 0 0 16 0 OUTPUT NODEFVAL "shiftout[15..0]"
-- Retrieval info: USED_PORT: taps0x 0 0 16 0 OUTPUT NODEFVAL "taps0x[15..0]"
-- Retrieval info: USED_PORT: taps100x 0 0 16 0 OUTPUT NODEFVAL "taps100x[15..0]"
-- Retrieval info: USED_PORT: taps101x 0 0 16 0 OUTPUT NODEFVAL "taps101x[15..0]"
-- Retrieval info: USED_PORT: taps102x 0 0 16 0 OUTPUT NODEFVAL "taps102x[15..0]"
-- Retrieval info: USED_PORT: taps103x 0 0 16 0 OUTPUT NODEFVAL "taps103x[15..0]"
-- Retrieval info: USED_PORT: taps104x 0 0 16 0 OUTPUT NODEFVAL "taps104x[15..0]"
-- Retrieval info: USED_PORT: taps105x 0 0 16 0 OUTPUT NODEFVAL "taps105x[15..0]"
-- Retrieval info: USED_PORT: taps106x 0 0 16 0 OUTPUT NODEFVAL "taps106x[15..0]"
-- Retrieval info: USED_PORT: taps107x 0 0 16 0 OUTPUT NODEFVAL "taps107x[15..0]"
-- Retrieval info: USED_PORT: taps108x 0 0 16 0 OUTPUT NODEFVAL "taps108x[15..0]"
-- Retrieval info: USED_PORT: taps109x 0 0 16 0 OUTPUT NODEFVAL "taps109x[15..0]"
-- Retrieval info: USED_PORT: taps10x 0 0 16 0 OUTPUT NODEFVAL "taps10x[15..0]"
-- Retrieval info: USED_PORT: taps110x 0 0 16 0 OUTPUT NODEFVAL "taps110x[15..0]"
-- Retrieval info: USED_PORT: taps111x 0 0 16 0 OUTPUT NODEFVAL "taps111x[15..0]"
-- Retrieval info: USED_PORT: taps112x 0 0 16 0 OUTPUT NODEFVAL "taps112x[15..0]"
-- Retrieval info: USED_PORT: taps113x 0 0 16 0 OUTPUT NODEFVAL "taps113x[15..0]"
-- Retrieval info: USED_PORT: taps114x 0 0 16 0 OUTPUT NODEFVAL "taps114x[15..0]"
-- Retrieval info: USED_PORT: taps115x 0 0 16 0 OUTPUT NODEFVAL "taps115x[15..0]"
-- Retrieval info: USED_PORT: taps116x 0 0 16 0 OUTPUT NODEFVAL "taps116x[15..0]"
-- Retrieval info: USED_PORT: taps117x 0 0 16 0 OUTPUT NODEFVAL "taps117x[15..0]"
-- Retrieval info: USED_PORT: taps118x 0 0 16 0 OUTPUT NODEFVAL "taps118x[15..0]"
-- Retrieval info: USED_PORT: taps119x 0 0 16 0 OUTPUT NODEFVAL "taps119x[15..0]"
-- Retrieval info: USED_PORT: taps11x 0 0 16 0 OUTPUT NODEFVAL "taps11x[15..0]"
-- Retrieval info: USED_PORT: taps120x 0 0 16 0 OUTPUT NODEFVAL "taps120x[15..0]"
-- Retrieval info: USED_PORT: taps121x 0 0 16 0 OUTPUT NODEFVAL "taps121x[15..0]"
-- Retrieval info: USED_PORT: taps122x 0 0 16 0 OUTPUT NODEFVAL "taps122x[15..0]"
-- Retrieval info: USED_PORT: taps123x 0 0 16 0 OUTPUT NODEFVAL "taps123x[15..0]"
-- Retrieval info: USED_PORT: taps124x 0 0 16 0 OUTPUT NODEFVAL "taps124x[15..0]"
-- Retrieval info: USED_PORT: taps125x 0 0 16 0 OUTPUT NODEFVAL "taps125x[15..0]"
-- Retrieval info: USED_PORT: taps126x 0 0 16 0 OUTPUT NODEFVAL "taps126x[15..0]"
-- Retrieval info: USED_PORT: taps127x 0 0 16 0 OUTPUT NODEFVAL "taps127x[15..0]"
-- Retrieval info: USED_PORT: taps12x 0 0 16 0 OUTPUT NODEFVAL "taps12x[15..0]"
-- Retrieval info: USED_PORT: taps13x 0 0 16 0 OUTPUT NODEFVAL "taps13x[15..0]"
-- Retrieval info: USED_PORT: taps14x 0 0 16 0 OUTPUT NODEFVAL "taps14x[15..0]"
-- Retrieval info: USED_PORT: taps15x 0 0 16 0 OUTPUT NODEFVAL "taps15x[15..0]"
-- Retrieval info: USED_PORT: taps16x 0 0 16 0 OUTPUT NODEFVAL "taps16x[15..0]"
-- Retrieval info: USED_PORT: taps17x 0 0 16 0 OUTPUT NODEFVAL "taps17x[15..0]"
-- Retrieval info: USED_PORT: taps18x 0 0 16 0 OUTPUT NODEFVAL "taps18x[15..0]"
-- Retrieval info: USED_PORT: taps19x 0 0 16 0 OUTPUT NODEFVAL "taps19x[15..0]"
-- Retrieval info: USED_PORT: taps1x 0 0 16 0 OUTPUT NODEFVAL "taps1x[15..0]"
-- Retrieval info: USED_PORT: taps20x 0 0 16 0 OUTPUT NODEFVAL "taps20x[15..0]"
-- Retrieval info: USED_PORT: taps21x 0 0 16 0 OUTPUT NODEFVAL "taps21x[15..0]"
-- Retrieval info: USED_PORT: taps22x 0 0 16 0 OUTPUT NODEFVAL "taps22x[15..0]"
-- Retrieval info: USED_PORT: taps23x 0 0 16 0 OUTPUT NODEFVAL "taps23x[15..0]"
-- Retrieval info: USED_PORT: taps24x 0 0 16 0 OUTPUT NODEFVAL "taps24x[15..0]"
-- Retrieval info: USED_PORT: taps25x 0 0 16 0 OUTPUT NODEFVAL "taps25x[15..0]"
-- Retrieval info: USED_PORT: taps26x 0 0 16 0 OUTPUT NODEFVAL "taps26x[15..0]"
-- Retrieval info: USED_PORT: taps27x 0 0 16 0 OUTPUT NODEFVAL "taps27x[15..0]"
-- Retrieval info: USED_PORT: taps28x 0 0 16 0 OUTPUT NODEFVAL "taps28x[15..0]"
-- Retrieval info: USED_PORT: taps29x 0 0 16 0 OUTPUT NODEFVAL "taps29x[15..0]"
-- Retrieval info: USED_PORT: taps2x 0 0 16 0 OUTPUT NODEFVAL "taps2x[15..0]"
-- Retrieval info: USED_PORT: taps30x 0 0 16 0 OUTPUT NODEFVAL "taps30x[15..0]"
-- Retrieval info: USED_PORT: taps31x 0 0 16 0 OUTPUT NODEFVAL "taps31x[15..0]"
-- Retrieval info: USED_PORT: taps32x 0 0 16 0 OUTPUT NODEFVAL "taps32x[15..0]"
-- Retrieval info: USED_PORT: taps33x 0 0 16 0 OUTPUT NODEFVAL "taps33x[15..0]"
-- Retrieval info: USED_PORT: taps34x 0 0 16 0 OUTPUT NODEFVAL "taps34x[15..0]"
-- Retrieval info: USED_PORT: taps35x 0 0 16 0 OUTPUT NODEFVAL "taps35x[15..0]"
-- Retrieval info: USED_PORT: taps36x 0 0 16 0 OUTPUT NODEFVAL "taps36x[15..0]"
-- Retrieval info: USED_PORT: taps37x 0 0 16 0 OUTPUT NODEFVAL "taps37x[15..0]"
-- Retrieval info: USED_PORT: taps38x 0 0 16 0 OUTPUT NODEFVAL "taps38x[15..0]"
-- Retrieval info: USED_PORT: taps39x 0 0 16 0 OUTPUT NODEFVAL "taps39x[15..0]"
-- Retrieval info: USED_PORT: taps3x 0 0 16 0 OUTPUT NODEFVAL "taps3x[15..0]"
-- Retrieval info: USED_PORT: taps40x 0 0 16 0 OUTPUT NODEFVAL "taps40x[15..0]"
-- Retrieval info: USED_PORT: taps41x 0 0 16 0 OUTPUT NODEFVAL "taps41x[15..0]"
-- Retrieval info: USED_PORT: taps42x 0 0 16 0 OUTPUT NODEFVAL "taps42x[15..0]"
-- Retrieval info: USED_PORT: taps43x 0 0 16 0 OUTPUT NODEFVAL "taps43x[15..0]"
-- Retrieval info: USED_PORT: taps44x 0 0 16 0 OUTPUT NODEFVAL "taps44x[15..0]"
-- Retrieval info: USED_PORT: taps45x 0 0 16 0 OUTPUT NODEFVAL "taps45x[15..0]"
-- Retrieval info: USED_PORT: taps46x 0 0 16 0 OUTPUT NODEFVAL "taps46x[15..0]"
-- Retrieval info: USED_PORT: taps47x 0 0 16 0 OUTPUT NODEFVAL "taps47x[15..0]"
-- Retrieval info: USED_PORT: taps48x 0 0 16 0 OUTPUT NODEFVAL "taps48x[15..0]"
-- Retrieval info: USED_PORT: taps49x 0 0 16 0 OUTPUT NODEFVAL "taps49x[15..0]"
-- Retrieval info: USED_PORT: taps4x 0 0 16 0 OUTPUT NODEFVAL "taps4x[15..0]"
-- Retrieval info: USED_PORT: taps50x 0 0 16 0 OUTPUT NODEFVAL "taps50x[15..0]"
-- Retrieval info: USED_PORT: taps51x 0 0 16 0 OUTPUT NODEFVAL "taps51x[15..0]"
-- Retrieval info: USED_PORT: taps52x 0 0 16 0 OUTPUT NODEFVAL "taps52x[15..0]"
-- Retrieval info: USED_PORT: taps53x 0 0 16 0 OUTPUT NODEFVAL "taps53x[15..0]"
-- Retrieval info: USED_PORT: taps54x 0 0 16 0 OUTPUT NODEFVAL "taps54x[15..0]"
-- Retrieval info: USED_PORT: taps55x 0 0 16 0 OUTPUT NODEFVAL "taps55x[15..0]"
-- Retrieval info: USED_PORT: taps56x 0 0 16 0 OUTPUT NODEFVAL "taps56x[15..0]"
-- Retrieval info: USED_PORT: taps57x 0 0 16 0 OUTPUT NODEFVAL "taps57x[15..0]"
-- Retrieval info: USED_PORT: taps58x 0 0 16 0 OUTPUT NODEFVAL "taps58x[15..0]"
-- Retrieval info: USED_PORT: taps59x 0 0 16 0 OUTPUT NODEFVAL "taps59x[15..0]"
-- Retrieval info: USED_PORT: taps5x 0 0 16 0 OUTPUT NODEFVAL "taps5x[15..0]"
-- Retrieval info: USED_PORT: taps60x 0 0 16 0 OUTPUT NODEFVAL "taps60x[15..0]"
-- Retrieval info: USED_PORT: taps61x 0 0 16 0 OUTPUT NODEFVAL "taps61x[15..0]"
-- Retrieval info: USED_PORT: taps62x 0 0 16 0 OUTPUT NODEFVAL "taps62x[15..0]"
-- Retrieval info: USED_PORT: taps63x 0 0 16 0 OUTPUT NODEFVAL "taps63x[15..0]"
-- Retrieval info: USED_PORT: taps64x 0 0 16 0 OUTPUT NODEFVAL "taps64x[15..0]"
-- Retrieval info: USED_PORT: taps65x 0 0 16 0 OUTPUT NODEFVAL "taps65x[15..0]"
-- Retrieval info: USED_PORT: taps66x 0 0 16 0 OUTPUT NODEFVAL "taps66x[15..0]"
-- Retrieval info: USED_PORT: taps67x 0 0 16 0 OUTPUT NODEFVAL "taps67x[15..0]"
-- Retrieval info: USED_PORT: taps68x 0 0 16 0 OUTPUT NODEFVAL "taps68x[15..0]"
-- Retrieval info: USED_PORT: taps69x 0 0 16 0 OUTPUT NODEFVAL "taps69x[15..0]"
-- Retrieval info: USED_PORT: taps6x 0 0 16 0 OUTPUT NODEFVAL "taps6x[15..0]"
-- Retrieval info: USED_PORT: taps70x 0 0 16 0 OUTPUT NODEFVAL "taps70x[15..0]"
-- Retrieval info: USED_PORT: taps71x 0 0 16 0 OUTPUT NODEFVAL "taps71x[15..0]"
-- Retrieval info: USED_PORT: taps72x 0 0 16 0 OUTPUT NODEFVAL "taps72x[15..0]"
-- Retrieval info: USED_PORT: taps73x 0 0 16 0 OUTPUT NODEFVAL "taps73x[15..0]"
-- Retrieval info: USED_PORT: taps74x 0 0 16 0 OUTPUT NODEFVAL "taps74x[15..0]"
-- Retrieval info: USED_PORT: taps75x 0 0 16 0 OUTPUT NODEFVAL "taps75x[15..0]"
-- Retrieval info: USED_PORT: taps76x 0 0 16 0 OUTPUT NODEFVAL "taps76x[15..0]"
-- Retrieval info: USED_PORT: taps77x 0 0 16 0 OUTPUT NODEFVAL "taps77x[15..0]"
-- Retrieval info: USED_PORT: taps78x 0 0 16 0 OUTPUT NODEFVAL "taps78x[15..0]"
-- Retrieval info: USED_PORT: taps79x 0 0 16 0 OUTPUT NODEFVAL "taps79x[15..0]"
-- Retrieval info: USED_PORT: taps7x 0 0 16 0 OUTPUT NODEFVAL "taps7x[15..0]"
-- Retrieval info: USED_PORT: taps80x 0 0 16 0 OUTPUT NODEFVAL "taps80x[15..0]"
-- Retrieval info: USED_PORT: taps81x 0 0 16 0 OUTPUT NODEFVAL "taps81x[15..0]"
-- Retrieval info: USED_PORT: taps82x 0 0 16 0 OUTPUT NODEFVAL "taps82x[15..0]"
-- Retrieval info: USED_PORT: taps83x 0 0 16 0 OUTPUT NODEFVAL "taps83x[15..0]"
-- Retrieval info: USED_PORT: taps84x 0 0 16 0 OUTPUT NODEFVAL "taps84x[15..0]"
-- Retrieval info: USED_PORT: taps85x 0 0 16 0 OUTPUT NODEFVAL "taps85x[15..0]"
-- Retrieval info: USED_PORT: taps86x 0 0 16 0 OUTPUT NODEFVAL "taps86x[15..0]"
-- Retrieval info: USED_PORT: taps87x 0 0 16 0 OUTPUT NODEFVAL "taps87x[15..0]"
-- Retrieval info: USED_PORT: taps88x 0 0 16 0 OUTPUT NODEFVAL "taps88x[15..0]"
-- Retrieval info: USED_PORT: taps89x 0 0 16 0 OUTPUT NODEFVAL "taps89x[15..0]"
-- Retrieval info: USED_PORT: taps8x 0 0 16 0 OUTPUT NODEFVAL "taps8x[15..0]"
-- Retrieval info: USED_PORT: taps90x 0 0 16 0 OUTPUT NODEFVAL "taps90x[15..0]"
-- Retrieval info: USED_PORT: taps91x 0 0 16 0 OUTPUT NODEFVAL "taps91x[15..0]"
-- Retrieval info: USED_PORT: taps92x 0 0 16 0 OUTPUT NODEFVAL "taps92x[15..0]"
-- Retrieval info: USED_PORT: taps93x 0 0 16 0 OUTPUT NODEFVAL "taps93x[15..0]"
-- Retrieval info: USED_PORT: taps94x 0 0 16 0 OUTPUT NODEFVAL "taps94x[15..0]"
-- Retrieval info: USED_PORT: taps95x 0 0 16 0 OUTPUT NODEFVAL "taps95x[15..0]"
-- Retrieval info: USED_PORT: taps96x 0 0 16 0 OUTPUT NODEFVAL "taps96x[15..0]"
-- Retrieval info: USED_PORT: taps97x 0 0 16 0 OUTPUT NODEFVAL "taps97x[15..0]"
-- Retrieval info: USED_PORT: taps98x 0 0 16 0 OUTPUT NODEFVAL "taps98x[15..0]"
-- Retrieval info: USED_PORT: taps99x 0 0 16 0 OUTPUT NODEFVAL "taps99x[15..0]"
-- Retrieval info: USED_PORT: taps9x 0 0 16 0 OUTPUT NODEFVAL "taps9x[15..0]"
-- Retrieval info: CONNECT: @clken 0 0 0 0 clken 0 0 0 0
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @shiftin 0 0 16 0 shiftin 0 0 16 0
-- Retrieval info: CONNECT: shiftout 0 0 16 0 @shiftout 0 0 16 0
-- Retrieval info: CONNECT: taps0x 0 0 16 0 @taps 0 0 16 0
-- Retrieval info: CONNECT: taps100x 0 0 16 0 @taps 0 0 16 1600
-- Retrieval info: CONNECT: taps101x 0 0 16 0 @taps 0 0 16 1616
-- Retrieval info: CONNECT: taps102x 0 0 16 0 @taps 0 0 16 1632
-- Retrieval info: CONNECT: taps103x 0 0 16 0 @taps 0 0 16 1648
-- Retrieval info: CONNECT: taps104x 0 0 16 0 @taps 0 0 16 1664
-- Retrieval info: CONNECT: taps105x 0 0 16 0 @taps 0 0 16 1680
-- Retrieval info: CONNECT: taps106x 0 0 16 0 @taps 0 0 16 1696
-- Retrieval info: CONNECT: taps107x 0 0 16 0 @taps 0 0 16 1712
-- Retrieval info: CONNECT: taps108x 0 0 16 0 @taps 0 0 16 1728
-- Retrieval info: CONNECT: taps109x 0 0 16 0 @taps 0 0 16 1744
-- Retrieval info: CONNECT: taps10x 0 0 16 0 @taps 0 0 16 160
-- Retrieval info: CONNECT: taps110x 0 0 16 0 @taps 0 0 16 1760
-- Retrieval info: CONNECT: taps111x 0 0 16 0 @taps 0 0 16 1776
-- Retrieval info: CONNECT: taps112x 0 0 16 0 @taps 0 0 16 1792
-- Retrieval info: CONNECT: taps113x 0 0 16 0 @taps 0 0 16 1808
-- Retrieval info: CONNECT: taps114x 0 0 16 0 @taps 0 0 16 1824
-- Retrieval info: CONNECT: taps115x 0 0 16 0 @taps 0 0 16 1840
-- Retrieval info: CONNECT: taps116x 0 0 16 0 @taps 0 0 16 1856
-- Retrieval info: CONNECT: taps117x 0 0 16 0 @taps 0 0 16 1872
-- Retrieval info: CONNECT: taps118x 0 0 16 0 @taps 0 0 16 1888
-- Retrieval info: CONNECT: taps119x 0 0 16 0 @taps 0 0 16 1904
-- Retrieval info: CONNECT: taps11x 0 0 16 0 @taps 0 0 16 176
-- Retrieval info: CONNECT: taps120x 0 0 16 0 @taps 0 0 16 1920
-- Retrieval info: CONNECT: taps121x 0 0 16 0 @taps 0 0 16 1936
-- Retrieval info: CONNECT: taps122x 0 0 16 0 @taps 0 0 16 1952
-- Retrieval info: CONNECT: taps123x 0 0 16 0 @taps 0 0 16 1968
-- Retrieval info: CONNECT: taps124x 0 0 16 0 @taps 0 0 16 1984
-- Retrieval info: CONNECT: taps125x 0 0 16 0 @taps 0 0 16 2000
-- Retrieval info: CONNECT: taps126x 0 0 16 0 @taps 0 0 16 2016
-- Retrieval info: CONNECT: taps127x 0 0 16 0 @taps 0 0 16 2032
-- Retrieval info: CONNECT: taps12x 0 0 16 0 @taps 0 0 16 192
-- Retrieval info: CONNECT: taps13x 0 0 16 0 @taps 0 0 16 208
-- Retrieval info: CONNECT: taps14x 0 0 16 0 @taps 0 0 16 224
-- Retrieval info: CONNECT: taps15x 0 0 16 0 @taps 0 0 16 240
-- Retrieval info: CONNECT: taps16x 0 0 16 0 @taps 0 0 16 256
-- Retrieval info: CONNECT: taps17x 0 0 16 0 @taps 0 0 16 272
-- Retrieval info: CONNECT: taps18x 0 0 16 0 @taps 0 0 16 288
-- Retrieval info: CONNECT: taps19x 0 0 16 0 @taps 0 0 16 304
-- Retrieval info: CONNECT: taps1x 0 0 16 0 @taps 0 0 16 16
-- Retrieval info: CONNECT: taps20x 0 0 16 0 @taps 0 0 16 320
-- Retrieval info: CONNECT: taps21x 0 0 16 0 @taps 0 0 16 336
-- Retrieval info: CONNECT: taps22x 0 0 16 0 @taps 0 0 16 352
-- Retrieval info: CONNECT: taps23x 0 0 16 0 @taps 0 0 16 368
-- Retrieval info: CONNECT: taps24x 0 0 16 0 @taps 0 0 16 384
-- Retrieval info: CONNECT: taps25x 0 0 16 0 @taps 0 0 16 400
-- Retrieval info: CONNECT: taps26x 0 0 16 0 @taps 0 0 16 416
-- Retrieval info: CONNECT: taps27x 0 0 16 0 @taps 0 0 16 432
-- Retrieval info: CONNECT: taps28x 0 0 16 0 @taps 0 0 16 448
-- Retrieval info: CONNECT: taps29x 0 0 16 0 @taps 0 0 16 464
-- Retrieval info: CONNECT: taps2x 0 0 16 0 @taps 0 0 16 32
-- Retrieval info: CONNECT: taps30x 0 0 16 0 @taps 0 0 16 480
-- Retrieval info: CONNECT: taps31x 0 0 16 0 @taps 0 0 16 496
-- Retrieval info: CONNECT: taps32x 0 0 16 0 @taps 0 0 16 512
-- Retrieval info: CONNECT: taps33x 0 0 16 0 @taps 0 0 16 528
-- Retrieval info: CONNECT: taps34x 0 0 16 0 @taps 0 0 16 544
-- Retrieval info: CONNECT: taps35x 0 0 16 0 @taps 0 0 16 560
-- Retrieval info: CONNECT: taps36x 0 0 16 0 @taps 0 0 16 576
-- Retrieval info: CONNECT: taps37x 0 0 16 0 @taps 0 0 16 592
-- Retrieval info: CONNECT: taps38x 0 0 16 0 @taps 0 0 16 608
-- Retrieval info: CONNECT: taps39x 0 0 16 0 @taps 0 0 16 624
-- Retrieval info: CONNECT: taps3x 0 0 16 0 @taps 0 0 16 48
-- Retrieval info: CONNECT: taps40x 0 0 16 0 @taps 0 0 16 640
-- Retrieval info: CONNECT: taps41x 0 0 16 0 @taps 0 0 16 656
-- Retrieval info: CONNECT: taps42x 0 0 16 0 @taps 0 0 16 672
-- Retrieval info: CONNECT: taps43x 0 0 16 0 @taps 0 0 16 688
-- Retrieval info: CONNECT: taps44x 0 0 16 0 @taps 0 0 16 704
-- Retrieval info: CONNECT: taps45x 0 0 16 0 @taps 0 0 16 720
-- Retrieval info: CONNECT: taps46x 0 0 16 0 @taps 0 0 16 736
-- Retrieval info: CONNECT: taps47x 0 0 16 0 @taps 0 0 16 752
-- Retrieval info: CONNECT: taps48x 0 0 16 0 @taps 0 0 16 768
-- Retrieval info: CONNECT: taps49x 0 0 16 0 @taps 0 0 16 784
-- Retrieval info: CONNECT: taps4x 0 0 16 0 @taps 0 0 16 64
-- Retrieval info: CONNECT: taps50x 0 0 16 0 @taps 0 0 16 800
-- Retrieval info: CONNECT: taps51x 0 0 16 0 @taps 0 0 16 816
-- Retrieval info: CONNECT: taps52x 0 0 16 0 @taps 0 0 16 832
-- Retrieval info: CONNECT: taps53x 0 0 16 0 @taps 0 0 16 848
-- Retrieval info: CONNECT: taps54x 0 0 16 0 @taps 0 0 16 864
-- Retrieval info: CONNECT: taps55x 0 0 16 0 @taps 0 0 16 880
-- Retrieval info: CONNECT: taps56x 0 0 16 0 @taps 0 0 16 896
-- Retrieval info: CONNECT: taps57x 0 0 16 0 @taps 0 0 16 912
-- Retrieval info: CONNECT: taps58x 0 0 16 0 @taps 0 0 16 928
-- Retrieval info: CONNECT: taps59x 0 0 16 0 @taps 0 0 16 944
-- Retrieval info: CONNECT: taps5x 0 0 16 0 @taps 0 0 16 80
-- Retrieval info: CONNECT: taps60x 0 0 16 0 @taps 0 0 16 960
-- Retrieval info: CONNECT: taps61x 0 0 16 0 @taps 0 0 16 976
-- Retrieval info: CONNECT: taps62x 0 0 16 0 @taps 0 0 16 992
-- Retrieval info: CONNECT: taps63x 0 0 16 0 @taps 0 0 16 1008
-- Retrieval info: CONNECT: taps64x 0 0 16 0 @taps 0 0 16 1024
-- Retrieval info: CONNECT: taps65x 0 0 16 0 @taps 0 0 16 1040
-- Retrieval info: CONNECT: taps66x 0 0 16 0 @taps 0 0 16 1056
-- Retrieval info: CONNECT: taps67x 0 0 16 0 @taps 0 0 16 1072
-- Retrieval info: CONNECT: taps68x 0 0 16 0 @taps 0 0 16 1088
-- Retrieval info: CONNECT: taps69x 0 0 16 0 @taps 0 0 16 1104
-- Retrieval info: CONNECT: taps6x 0 0 16 0 @taps 0 0 16 96
-- Retrieval info: CONNECT: taps70x 0 0 16 0 @taps 0 0 16 1120
-- Retrieval info: CONNECT: taps71x 0 0 16 0 @taps 0 0 16 1136
-- Retrieval info: CONNECT: taps72x 0 0 16 0 @taps 0 0 16 1152
-- Retrieval info: CONNECT: taps73x 0 0 16 0 @taps 0 0 16 1168
-- Retrieval info: CONNECT: taps74x 0 0 16 0 @taps 0 0 16 1184
-- Retrieval info: CONNECT: taps75x 0 0 16 0 @taps 0 0 16 1200
-- Retrieval info: CONNECT: taps76x 0 0 16 0 @taps 0 0 16 1216
-- Retrieval info: CONNECT: taps77x 0 0 16 0 @taps 0 0 16 1232
-- Retrieval info: CONNECT: taps78x 0 0 16 0 @taps 0 0 16 1248
-- Retrieval info: CONNECT: taps79x 0 0 16 0 @taps 0 0 16 1264
-- Retrieval info: CONNECT: taps7x 0 0 16 0 @taps 0 0 16 112
-- Retrieval info: CONNECT: taps80x 0 0 16 0 @taps 0 0 16 1280
-- Retrieval info: CONNECT: taps81x 0 0 16 0 @taps 0 0 16 1296
-- Retrieval info: CONNECT: taps82x 0 0 16 0 @taps 0 0 16 1312
-- Retrieval info: CONNECT: taps83x 0 0 16 0 @taps 0 0 16 1328
-- Retrieval info: CONNECT: taps84x 0 0 16 0 @taps 0 0 16 1344
-- Retrieval info: CONNECT: taps85x 0 0 16 0 @taps 0 0 16 1360
-- Retrieval info: CONNECT: taps86x 0 0 16 0 @taps 0 0 16 1376
-- Retrieval info: CONNECT: taps87x 0 0 16 0 @taps 0 0 16 1392
-- Retrieval info: CONNECT: taps88x 0 0 16 0 @taps 0 0 16 1408
-- Retrieval info: CONNECT: taps89x 0 0 16 0 @taps 0 0 16 1424
-- Retrieval info: CONNECT: taps8x 0 0 16 0 @taps 0 0 16 128
-- Retrieval info: CONNECT: taps90x 0 0 16 0 @taps 0 0 16 1440
-- Retrieval info: CONNECT: taps91x 0 0 16 0 @taps 0 0 16 1456
-- Retrieval info: CONNECT: taps92x 0 0 16 0 @taps 0 0 16 1472
-- Retrieval info: CONNECT: taps93x 0 0 16 0 @taps 0 0 16 1488
-- Retrieval info: CONNECT: taps94x 0 0 16 0 @taps 0 0 16 1504
-- Retrieval info: CONNECT: taps95x 0 0 16 0 @taps 0 0 16 1520
-- Retrieval info: CONNECT: taps96x 0 0 16 0 @taps 0 0 16 1536
-- Retrieval info: CONNECT: taps97x 0 0 16 0 @taps 0 0 16 1552
-- Retrieval info: CONNECT: taps98x 0 0 16 0 @taps 0 0 16 1568
-- Retrieval info: CONNECT: taps99x 0 0 16 0 @taps 0 0 16 1584
-- Retrieval info: CONNECT: taps9x 0 0 16 0 @taps 0 0 16 144
-- Retrieval info: GEN_FILE: TYPE_NORMAL Shift_registers_128.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Shift_registers_128.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Shift_registers_128.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Shift_registers_128.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Shift_registers_128_inst.vhd TRUE
-- Retrieval info: LIB_FILE: altera_mf
