library IEEE;
use IEEE.STD_LOGIC_1164.ALL;  
use IEEE.NUMERIC_STD.ALL;
use work.data_types.all;

entity impulsebench is
end;

architecture testbench of impulsebench is

	signal rst : std_logic := '0';
	signal clk : std_logic := '0';
	signal interclk : std_logic := '0';
	signal sndclk : std_logic := '0';
	signal word : signed(0 downto 0);
	signal inter : signed(15 downto 0);
  signal resp : signed(15 downto 0);

  component polyphase
    Generic (
        coef_scale : integer := 1024;
        w_acc : integer := 32;
        w_in : integer := 16;
        w_out : integer := 16;
        coef : array_of_integers := (1, -5, -17, -24, 3, 83, 194, 277, 277, 194, 83, 3, -24, -17, -5, 1);
        D : integer := 4
    );
    port (
      rst    : in std_logic;
      clk    : in std_logic;
      inclk : in std_logic;
      outclk : out std_logic;
      word   : in signed(w_in-1 downto 0);
      resp   : out signed(w_out-1 downto 0)
    );
  end component;

    
begin
  rst <= '1' AFTER 20 ns; -- reset pin
  clk <= NOT clk AFTER 10 ns; -- "fast clock"; 50 MHz klok

  process(clk)
    variable counter: integer := 0;
  begin
    if rising_edge(clk) then
      counter := counter + 1;
      if counter < 3000 then
        word <= "0";
      elsif counter < 100000 then
        word <= "1";
      else
        word <= not word;
      end if;
    end if;
  end process;

  filter_inst1 : polyphase
  generic map (
    coef_scale => 1,
    w_acc => 32,
    w_in => 1,
    w_out => 16,
    D => 64,
    coef => (
-2,-2,-5,-9,-13,-16,-16,-10,4,26,58,98,140,182,216,239,246,237,213,177,135,92,54,23,2,-11,-16,-16,-12,-8,-5,-2,
-1,-3,-5,-9,-13,-16,-15,-9,6,30,63,103,146,187,220,241,246,235,209,172,130,87,50,20,-1,-12,-16,-15,-12,-8,-4,-2,
-1,-3,-6,-10,-14,-16,-15,-7,8,34,68,108,151,191,223,242,245,232,204,167,124,82,45,17,-2,-13,-16,-15,-11,-7,-4,-2,
-1,-3,-6,-10,-14,-16,-14,-6,11,37,72,113,156,196,226,243,244,229,200,162,119,77,41,14,-4,-14,-16,-15,-11,-7,-3,-1,
-1,-3,-7,-11,-15,-16,-14,-4,14,41,77,119,162,200,229,244,243,226,196,156,113,72,37,11,-6,-14,-16,-14,-10,-6,-3,-1,
-2,-4,-7,-11,-15,-16,-13,-2,17,45,82,124,167,204,232,245,242,223,191,151,108,68,34,8,-7,-15,-16,-14,-10,-6,-3,-1,
-2,-4,-8,-12,-15,-16,-12,-1,20,50,87,130,172,209,235,246,241,220,187,146,103,63,30,6,-9,-15,-16,-13,-9,-5,-3,-1,
-2,-5,-8,-12,-16,-16,-11,2,23,54,92,135,177,213,237,246,239,216,182,140,98,58,26,4,-10,-16,-16,-13,-9,-5,-2,-2
  )
  )
  port map (
    rst => rst,
    clk => clk,
    inclk => clk,
    outclk => interclk,
    word => word,
    resp => inter
  );
  filter_inst2 : polyphase
  generic map (
    coef_scale => 2**16,
    w_acc => 32,
    w_in => 16,
    w_out => 16,
    D => 16,
    coef => (
34,-9,12,-17,20,-18,8,12,-44,88,-145,211,-282,354,-428,531,3672,289,-326,306,-262,209,-152,100,-56,23,-1,-11,16,-15,11,-9,
0,-9,13,-19,23,-24,18,-1,-29,73,-133,207,-293,393,-522,790,3634,67,-221,250,-235,200,-155,109,-67,34,-10,-5,11,-13,10,-9,
0,-8,13,-20,26,-30,27,-14,-13,56,-116,196,-296,422,-607,1060,3559,-133,-116,190,-202,185,-152,113,-75,43,-18,2,7,-10,9,-8,
-0,-8,12,-21,29,-35,35,-27,4,35,-95,178,-289,439,-678,1339,3447,-308,-14,126,-165,165,-145,114,-81,50,-26,8,2,-7,7,-8,
-1,-7,12,-21,30,-39,43,-39,22,13,-70,155,-273,443,-733,1621,3301,-456,82,61,-123,141,-134,112,-84,56,-32,14,-2,-4,5,-7,
-1,-5,10,-20,31,-42,50,-51,39,-10,-43,125,-247,433,-769,1902,3125,-577,171,-2,-79,114,-119,106,-84,60,-37,19,-6,-1,3,-6,
-2,-4,9,-18,30,-44,55,-61,56,-34,-12,90,-212,408,-782,2178,2920,-670,249,-63,-35,83,-100,97,-82,62,-41,23,-10,2,1,-5,
-3,-2,7,-16,29,-44,59,-70,72,-57,19,51,-169,369,-771,2442,2691,-734,315,-119,9,52,-80,86,-77,61,-43,26,-13,4,-0,-4,
-4,-0,4,-13,26,-43,61,-77,86,-80,52,9,-119,315,-734,2691,2442,-771,369,-169,51,19,-57,72,-70,59,-44,29,-16,7,-2,-3,
-5,1,2,-10,23,-41,62,-82,97,-100,83,-35,-63,249,-670,2920,2178,-782,408,-212,90,-12,-34,56,-61,55,-44,30,-18,9,-4,-2,
-6,3,-1,-6,19,-37,60,-84,106,-119,114,-79,-2,171,-577,3125,1902,-769,433,-247,125,-43,-10,39,-51,50,-42,31,-20,10,-5,-1,
-7,5,-4,-2,14,-32,56,-84,112,-134,141,-123,61,82,-456,3301,1621,-733,443,-273,155,-70,13,22,-39,43,-39,30,-21,12,-7,-1,
-8,7,-7,2,8,-26,50,-81,114,-145,165,-165,126,-14,-308,3447,1339,-678,439,-289,178,-95,35,4,-27,35,-35,29,-21,12,-8,-0,
-8,9,-10,7,2,-18,43,-75,113,-152,185,-202,190,-116,-133,3559,1060,-607,422,-296,196,-116,56,-13,-14,27,-30,26,-20,13,-8,0,
-9,10,-13,11,-5,-10,34,-67,109,-155,200,-235,250,-221,67,3634,790,-522,393,-293,207,-133,73,-29,-1,18,-24,23,-19,13,-9,0,
-9,11,-15,16,-11,-1,23,-56,100,-152,209,-262,306,-326,289,3672,531,-428,354,-282,211,-145,88,-44,12,8,-18,20,-17,12,-9,34
  )
  )
  port map (
    rst => rst,
    clk => clk,
    inclk => interclk,
    outclk => sndclk,
    word => inter,
    resp => resp
  );
end;
