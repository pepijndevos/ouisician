library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity WahWah_FX is
port (
	CLK_50		: in std_logic;
	nReset		: in std_logic;
	new_val		: in std_logic;       -- indicates a new input value, input from data_over
	data_in		: in signed (15 downto 0);         
	data_out		: out signed (15 downto 0);   -- Output
	filterid: IN std_logic_vector(7 DOWNTO 0);
	chan: IN std_logic_vector(7 DOWNTO 0);
	fil_data: IN std_logic_vector(31 DOWNTO 0)
);
end entity WahWah_FX;

architecture behaviour of WahWah_FX is
constant W_coef : integer := 23;
constant W_in : integer := 16;
constant A0 : integer :=1048576 ;
constant A2 : integer :=982099 ;
constant B0 : integer :=33239 ;
constant B1 : integer := 0;
constant B2 : integer := -33239 ; 
constant Arr_size : integer := 3456;

component IIRDF1_BW is
generic (
   W_in : integer ;
	W_coef : integer;
	A0 : integer;
	A2 : integer;
	B0 : integer;
	B1 : integer;
	B2 : integer    
);
port (
	iCLK            : in std_logic;
	iRESET_N        : in std_logic;
	new_val         : in std_logic;       -- indicates a new input value, input from data_over
	IIR_in          : in signed (15 downto 0);   -- singed is expected             
	IIR_out         : out signed (15 downto 0);   -- Output
   A1 : in signed(W_coef-1 downto 0)

);
end component;


type cA1_array_type is array (0 to Arr_size) of integer;
signal A1 : cA1_array_type:=(-2029624,-2029618,-2029611,-2029605,-2029599,-2029592,-2029586,-2029579,-2029573,-2029567,-2029560,-2029554,-2029547,-2029541,-2029534,-2029528,-2029521,-2029515,-2029508,-2029502,-2029495,-2029489,-2029482,-2029475,-2029469,-2029462,-2029456,-2029449,-2029443,-2029436,-2029429,-2029423,-2029416,-2029409,-2029403,-2029396,-2029389,-2029383,-2029376,-2029369,-2029362,-2029356,-2029349,-2029342,-2029335,-2029329,-2029322,-2029315,-2029308,-2029301,-2029295,-2029288,-2029281,-2029274,-2029267,-2029260,-2029254,-2029247,-2029240,-2029233,-2029226,-2029219,-2029212,-2029205,-2029198,-2029191,-2029184,-2029177,-2029170,-2029163,-2029156,-2029149,-2029142,-2029135,-2029128,-2029121,-2029114,-2029107,-2029100,-2029093,-2029086,-2029079,-2029071,-2029064,-2029057,-2029050,-2029043,-2029036,-2029028,-2029021,-2029014,-2029007,-2029000,-2028992,-2028985,-2028978,-2028971,-2028963,-2028956,-2028949,-2028942,-2028934,-2028927,-2028920,-2028912,-2028905,-2028898,-2028890,-2028883,-2028876,-2028868,-2028861,-2028853,-2028846,-2028839,-2028831,-2028824,-2028816,-2028809,-2028801,-2028794,-2028786,-2028779,-2028771,-2028764,-2028756,-2028749,-2028741,-2028734,-2028726,-2028718,-2028711,-2028703,-2028696,-2028688,-2028680,-2028673,-2028665,-2028658,-2028650,-2028642,-2028635,-2028627,-2028619,-2028611,-2028604,-2028596,-2028588,-2028580,-2028573,-2028565,-2028557,-2028549,-2028542,-2028534,-2028526,-2028518,-2028510,-2028503,-2028495,-2028487,-2028479,-2028471,-2028463,-2028455,-2028447,-2028439,-2028432,-2028424,-2028416,-2028408,-2028400,-2028392,-2028384,-2028376,-2028368,-2028360,-2028352,-2028344,-2028336,-2028328,-2028320,-2028312,-2028303,-2028295,-2028287,-2028279,-2028271,-2028263,-2028255,-2028247,-2028239,-2028230,-2028222,-2028214,-2028206,-2028198,-2028189,-2028181,-2028173,-2028165,-2028157,-2028148,-2028140,-2028132,-2028123,-2028115,-2028107,-2028099,-2028090,-2028082,-2028074,-2028065,-2028057,-2028049,-2028040,-2028032,-2028023,-2028015,-2028007,-2027998,-2027990,-2027981,-2027973,-2027964,-2027956,-2027947,-2027939,-2027930,-2027922,-2027913,-2027905,-2027896,-2027888,-2027879,-2027871,-2027862,-2027853,-2027845,-2027836,-2027828,-2027819,-2027810,-2027802,-2027793,-2027784,-2027776,-2027767,-2027758,-2027750,-2027741,-2027732,-2027724,-2027715,-2027706,-2027697,-2027689,-2027680,-2027671,-2027662,-2027653,-2027645,-2027636,-2027627,-2027618,-2027609,-2027600,-2027592,-2027583,-2027574,-2027565,-2027556,-2027547,-2027538,-2027529,-2027520,-2027511,-2027502,-2027493,-2027484,-2027475,-2027466,-2027457,-2027448,-2027439,-2027430,-2027421,-2027412,-2027403,-2027394,-2027385,-2027376,-2027367,-2027358,-2027349,-2027339,-2027330,-2027321,-2027312,-2027303,-2027294,-2027285,-2027275,-2027266,-2027257,-2027248,-2027238,-2027229,-2027220,-2027211,-2027201,-2027192,-2027183,-2027174,-2027164,-2027155,-2027146,-2027136,-2027127,-2027118,-2027108,-2027099,-2027089,-2027080,-2027071,-2027061,-2027052,-2027042,-2027033,-2027023,-2027014,-2027005,-2026995,-2026986,-2026976,-2026967,-2026957,-2026948,-2026938,-2026928,-2026919,-2026909,-2026900,-2026890,-2026881,-2026871,-2026861,-2026852,-2026842,-2026832,-2026823,-2026813,-2026803,-2026794,-2026784,-2026774,-2026765,-2026755,-2026745,-2026736,-2026726,-2026716,-2026706,-2026697,-2026687,-2026677,-2026667,-2026657,-2026648,-2026638,-2026628,-2026618,-2026608,-2026598,-2026588,-2026579,-2026569,-2026559,-2026549,-2026539,-2026529,-2026519,-2026509,-2026499,-2026489,-2026479,-2026469,-2026459,-2026449,-2026439,-2026429,-2026419,-2026409,-2026399,-2026389,-2026379,-2026369,-2026359,-2026349,-2026338,-2026328,-2026318,-2026308,-2026298,-2026288,-2026278,-2026267,-2026257,-2026247,-2026237,-2026227,-2026216,-2026206,-2026196,-2026186,-2026175,-2026165,-2026155,-2026145,-2026134,-2026124,-2026114,-2026103,-2026093,-2026083,-2026072,-2026062,-2026052,-2026041,-2026031,-2026020,-2026010,-2026000,-2025989,-2025979,-2025968,-2025958,-2025947,-2025937,-2025926,-2025916,-2025905,-2025895,-2025884,-2025874,-2025863,-2025853,-2025842,-2025832,-2025821,-2025810,-2025800,-2025789,-2025779,-2025768,-2025757,-2025747,-2025736,-2025725,-2025715,-2025704,-2025693,-2025683,-2025672,-2025661,-2025650,-2025640,-2025629,-2025618,-2025607,-2025597,-2025586,-2025575,-2025564,-2025553,-2025543,-2025532,-2025521,-2025510,-2025499,-2025488,-2025477,-2025467,-2025456,-2025445,-2025434,-2025423,-2025412,-2025401,-2025390,-2025379,-2025368,-2025357,-2025346,-2025335,-2025324,-2025313,-2025302,-2025291,-2025280,-2025269,-2025258,-2025247,-2025236,-2025225,-2025213,-2025202,-2025191,-2025180,-2025169,-2025158,-2025147,-2025135,-2025124,-2025113,-2025102,-2025091,-2025079,-2025068,-2025057,-2025046,-2025034,-2025023,-2025012,-2025001,-2024989,-2024978,-2024967,-2024955,-2024944,-2024933,-2024921,-2024910,-2024899,-2024887,-2024876,-2024864,-2024853,-2024842,-2024830,-2024819,-2024807,-2024796,-2024784,-2024773,-2024761,-2024750,-2024738,-2024727,-2024715,-2024704,-2024692,-2024681,-2024669,-2024658,-2024646,-2024634,-2024623,-2024611,-2024600,-2024588,-2024576,-2024565,-2024553,-2024541,-2024530,-2024518,-2024506,-2024495,-2024483,-2024471,-2024459,-2024448,-2024436,-2024424,-2024412,-2024401,-2024389,-2024377,-2024365,-2024353,-2024342,-2024330,-2024318,-2024306,-2024294,-2024282,-2024271,-2024259,-2024247,-2024235,-2024223,-2024211,-2024199,-2024187,-2024175,-2024163,-2024151,-2024139,-2024127,-2024115,-2024103,-2024091,-2024079,-2024067,-2024055,-2024043,-2024031,-2024019,-2024007,-2023995,-2023983,-2023970,-2023958,-2023946,-2023934,-2023922,-2023910,-2023898,-2023885,-2023873,-2023861,-2023849,-2023837,-2023824,-2023812,-2023800,-2023788,-2023775,-2023763,-2023751,-2023739,-2023726,-2023714,-2023702,-2023689,-2023677,-2023665,-2023652,-2023640,-2023627,-2023615,-2023603,-2023590,-2023578,-2023565,-2023553,-2023541,-2023528,-2023516,-2023503,-2023491,-2023478,-2023466,-2023453,-2023441,-2023428,-2023416,-2023403,-2023390,-2023378,-2023365,-2023353,-2023340,-2023328,-2023315,-2023302,-2023290,-2023277,-2023264,-2023252,-2023239,-2023226,-2023214,-2023201,-2023188,-2023176,-2023163,-2023150,-2023137,-2023125,-2023112,-2023099,-2023086,-2023073,-2023061,-2023048,-2023035,-2023022,-2023009,-2022997,-2022984,-2022971,-2022958,-2022945,-2022932,-2022919,-2022906,-2022893,-2022880,-2022868,-2022855,-2022842,-2022829,-2022816,-2022803,-2022790,-2022777,-2022764,-2022751,-2022738,-2022725,-2022711,-2022698,-2022685,-2022672,-2022659,-2022646,-2022633,-2022620,-2022607,-2022594,-2022580,-2022567,-2022554,-2022541,-2022528,-2022515,-2022501,-2022488,-2022475,-2022462,-2022448,-2022435,-2022422,-2022409,-2022395,-2022382,-2022369,-2022355,-2022342,-2022329,-2022315,-2022302,-2022289,-2022275,-2022262,-2022249,-2022235,-2022222,-2022208,-2022195,-2022182,-2022168,-2022155,-2022141,-2022128,-2022114,-2022101,-2022087,-2022074,-2022060,-2022047,-2022033,-2022020,-2022006,-2021993,-2021979,-2021965,-2021952,-2021938,-2021925,-2021911,-2021897,-2021884,-2021870,-2021856,-2021843,-2021829,-2021815,-2021802,-2021788,-2021774,-2021760,-2021747,-2021733,-2021719,-2021706,-2021692,-2021678,-2021664,-2021650,-2021637,-2021623,-2021609,-2021595,-2021581,-2021567,-2021554,-2021540,-2021526,-2021512,-2021498,-2021484,-2021470,-2021456,-2021442,-2021428,-2021414,-2021400,-2021386,-2021372,-2021358,-2021344,-2021330,-2021316,-2021302,-2021288,-2021274,-2021260,-2021246,-2021232,-2021218,-2021204,-2021190,-2021176,-2021162,-2021147,-2021133,-2021119,-2021105,-2021091,-2021077,-2021062,-2021048,-2021034,-2021020,-2021006,-2020991,-2020977,-2020963,-2020948,-2020934,-2020920,-2020906,-2020891,-2020877,-2020863,-2020848,-2020834,-2020820,-2020805,-2020791,-2020777,-2020762,-2020748,-2020733,-2020719,-2020704,-2020690,-2020676,-2020661,-2020647,-2020632,-2020618,-2020603,-2020589,-2020574,-2020560,-2020545,-2020531,-2020516,-2020502,-2020487,-2020472,-2020458,-2020443,-2020429,-2020414,-2020399,-2020385,-2020370,-2020355,-2020341,-2020326,-2020311,-2020297,-2020282,-2020267,-2020253,-2020238,-2020223,-2020208,-2020194,-2020179,-2020164,-2020149,-2020134,-2020120,-2020105,-2020090,-2020075,-2020060,-2020046,-2020031,-2020016,-2020001,-2019986,-2019971,-2019956,-2019941,-2019926,-2019911,-2019897,-2019882,-2019867,-2019852,-2019837,-2019822,-2019807,-2019792,-2019777,-2019762,-2019747,-2019732,-2019716,-2019701,-2019686,-2019671,-2019656,-2019641,-2019626,-2019611,-2019596,-2019581,-2019565,-2019550,-2019535,-2019520,-2019505,-2019489,-2019474,-2019459,-2019444,-2019429,-2019413,-2019398,-2019383,-2019368,-2019352,-2019337,-2019322,-2019306,-2019291,-2019276,-2019260,-2019245,-2019230,-2019214,-2019199,-2019184,-2019168,-2019153,-2019137,-2019122,-2019106,-2019091,-2019076,-2019060,-2019045,-2019029,-2019014,-2018998,-2018983,-2018967,-2018952,-2018936,-2018921,-2018905,-2018889,-2018874,-2018858,-2018843,-2018827,-2018812,-2018796,-2018780,-2018765,-2018749,-2018733,-2018718,-2018702,-2018686,-2018671,-2018655,-2018639,-2018623,-2018608,-2018592,-2018576,-2018560,-2018545,-2018529,-2018513,-2018497,-2018482,-2018466,-2018450,-2018434,-2018418,-2018402,-2018386,-2018371,-2018355,-2018339,-2018323,-2018307,-2018291,-2018275,-2018259,-2018243,-2018227,-2018211,-2018195,-2018179,-2018163,-2018147,-2018131,-2018115,-2018099,-2018083,-2018067,-2018051,-2018035,-2018019,-2018003,-2017987,-2017971,-2017955,-2017938,-2017922,-2017906,-2017890,-2017874,-2017858,-2017842,-2017825,-2017809,-2017793,-2017777,-2017760,-2017744,-2017728,-2017712,-2017695,-2017679,-2017663,-2017647,-2017630,-2017614,-2017598,-2017581,-2017565,-2017549,-2017532,-2017516,-2017500,-2017483,-2017467,-2017450,-2017434,-2017417,-2017401,-2017385,-2017368,-2017352,-2017335,-2017319,-2017302,-2017286,-2017269,-2017253,-2017236,-2017220,-2017203,-2017187,-2017170,-2017153,-2017137,-2017120,-2017104,-2017087,-2017070,-2017054,-2017037,-2017020,-2017004,-2016987,-2016970,-2016954,-2016937,-2016920,-2016904,-2016887,-2016870,-2016853,-2016837,-2016820,-2016803,-2016786,-2016770,-2016753,-2016736,-2016719,-2016702,-2016685,-2016669,-2016652,-2016635,-2016618,-2016601,-2016584,-2016567,-2016550,-2016533,-2016517,-2016500,-2016483,-2016466,-2016449,-2016432,-2016415,-2016398,-2016381,-2016364,-2016347,-2016330,-2016313,-2016296,-2016278,-2016261,-2016244,-2016227,-2016210,-2016193,-2016176,-2016159,-2016142,-2016124,-2016107,-2016090,-2016073,-2016056,-2016039,-2016021,-2016004,-2015987,-2015970,-2015952,-2015935,-2015918,-2015901,-2015883,-2015866,-2015849,-2015832,-2015814,-2015797,-2015780,-2015762,-2015745,-2015727,-2015710,-2015693,-2015675,-2015658,-2015641,-2015623,-2015606,-2015588,-2015571,-2015553,-2015536,-2015518,-2015501,-2015483,-2015466,-2015448,-2015431,-2015413,-2015396,-2015378,-2015361,-2015343,-2015326,-2015308,-2015290,-2015273,-2015255,-2015237,-2015220,-2015202,-2015185,-2015167,-2015149,-2015132,-2015114,-2015096,-2015078,-2015061,-2015043,-2015025,-2015007,-2014990,-2014972,-2014954,-2014936,-2014919,-2014901,-2014883,-2014865,-2014847,-2014830,-2014812,-2014794,-2014776,-2014758,-2014740,-2014722,-2014704,-2014686,-2014669,-2014651,-2014633,-2014615,-2014597,-2014579,-2014561,-2014543,-2014525,-2014507,-2014489,-2014471,-2014453,-2014435,-2014417,-2014398,-2014380,-2014362,-2014344,-2014326,-2014308,-2014290,-2014272,-2014254,-2014235,-2014217,-2014199,-2014181,-2014163,-2014145,-2014126,-2014108,-2014090,-2014072,-2014053,-2014035,-2014017,-2013999,-2013980,-2013962,-2013944,-2013925,-2013907,-2013889,-2013870,-2013852,-2013834,-2013815,-2013797,-2013779,-2013760,-2013742,-2013723,-2013705,-2013687,-2013668,-2013650,-2013631,-2013613,-2013594,-2013576,-2013557,-2013539,-2013520,-2013502,-2013483,-2013465,-2013446,-2013428,-2013409,-2013390,-2013372,-2013353,-2013335,-2013316,-2013297,-2013279,-2013260,-2013241,-2013223,-2013204,-2013185,-2013167,-2013148,-2013129,-2013111,-2013092,-2013073,-2013054,-2013036,-2013017,-2012998,-2012979,-2012960,-2012942,-2012923,-2012904,-2012885,-2012866,-2012848,-2012829,-2012810,-2012791,-2012772,-2012753,-2012734,-2012715,-2012696,-2012677,-2012658,-2012640,-2012621,-2012602,-2012583,-2012564,-2012545,-2012526,-2012507,-2012488,-2012468,-2012449,-2012430,-2012411,-2012392,-2012373,-2012354,-2012335,-2012316,-2012297,-2012278,-2012258,-2012239,-2012220,-2012201,-2012182,-2012163,-2012143,-2012124,-2012105,-2012086,-2012066,-2012047,-2012028,-2012009,-2011989,-2011970,-2011951,-2011932,-2011912,-2011893,-2011874,-2011854,-2011835,-2011816,-2011796,-2011777,-2011757,-2011738,-2011719,-2011699,-2011680,-2011660,-2011641,-2011621,-2011602,-2011583,-2011563,-2011544,-2011524,-2011505,-2011485,-2011466,-2011446,-2011426,-2011407,-2011387,-2011368,-2011348,-2011329,-2011309,-2011289,-2011270,-2011250,-2011230,-2011211,-2011191,-2011172,-2011152,-2011132,-2011112,-2011093,-2011073,-2011053,-2011034,-2011014,-2010994,-2010974,-2010955,-2010935,-2010915,-2010895,-2010875,-2010856,-2010836,-2010816,-2010796,-2010776,-2010756,-2010737,-2010717,-2010697,-2010677,-2010657,-2010637,-2010617,-2010597,-2010577,-2010557,-2010537,-2010517,-2010497,-2010477,-2010457,-2010437,-2010417,-2010397,-2010377,-2010357,-2010337,-2010317,-2010297,-2010277,-2010257,-2010237,-2010217,-2010196,-2010176,-2010156,-2010136,-2010116,-2010096,-2010075,-2010055,-2010035,-2010015,-2009995,-2009974,-2009954,-2009934,-2009914,-2009893,-2009873,-2009853,-2009833,-2009812,-2009792,-2009772,-2009751,-2009731,-2009711,-2009690,-2009670,-2009650,-2009629,-2009609,-2009588,-2009568,-2009548,-2009527,-2009507,-2009486,-2009466,-2009445,-2009425,-2009404,-2009384,-2009363,-2009343,-2009322,-2009302,-2009281,-2009261,-2009240,-2009219,-2009199,-2009178,-2009158,-2009137,-2009116,-2009096,-2009075,-2009055,-2009034,-2009013,-2008993,-2008972,-2008951,-2008930,-2008910,-2008889,-2008868,-2008848,-2008827,-2008806,-2008785,-2008765,-2008744,-2008723,-2008702,-2008681,-2008660,-2008640,-2008619,-2008598,-2008577,-2008556,-2008535,-2008514,-2008494,-2008473,-2008452,-2008431,-2008410,-2008389,-2008368,-2008347,-2008326,-2008305,-2008284,-2008263,-2008242,-2008221,-2008200,-2008179,-2008158,-2008137,-2008116,-2008095,-2008074,-2008053,-2008031,-2008010,-2007989,-2007968,-2007947,-2007926,-2007905,-2007883,-2007862,-2007841,-2007820,-2007799,-2007777,-2007756,-2007735,-2007714,-2007692,-2007671,-2007650,-2007629,-2007607,-2007586,-2007565,-2007543,-2007522,-2007501,-2007479,-2007458,-2007437,-2007415,-2007394,-2007373,-2007351,-2007330,-2007308,-2007287,-2007265,-2007244,-2007223,-2007201,-2007180,-2007158,-2007137,-2007115,-2007094,-2007072,-2007051,-2007029,-2007007,-2006986,-2006964,-2006943,-2006921,-2006900,-2006878,-2006856,-2006835,-2006813,-2006791,-2006770,-2006748,-2006726,-2006705,-2006683,-2006661,-2006640,-2006618,-2006596,-2006574,-2006553,-2006531,-2006509,-2006487,-2006466,-2006444,-2006422,-2006400,-2006378,-2006357,-2006335,-2006313,-2006291,-2006269,-2006247,-2006225,-2006203,-2006182,-2006160,-2006138,-2006116,-2006094,-2006072,-2006050,-2006028,-2006006,-2005984,-2005962,-2005940,-2005918,-2005896,-2005874,-2005852,-2005830,-2005808,-2005786,-2005764,-2005741,-2005719,-2005697,-2005675,-2005653,-2005631,-2005609,-2005586,-2005564,-2005542,-2005520,-2005498,-2005476,-2005453,-2005431,-2005409,-2005387,-2005364,-2005342,-2005320,-2005298,-2005275,-2005253,-2005231,-2005208,-2005186,-2005164,-2005141,-2005119,-2005097,-2005074,-2005052,-2005029,-2005007,-2004985,-2004962,-2004940,-2004917,-2004895,-2004872,-2004850,-2004828,-2004805,-2004783,-2004760,-2004738,-2004715,-2004693,-2004670,-2004647,-2004625,-2004602,-2004580,-2004557,-2004535,-2004512,-2004489,-2004467,-2004444,-2004421,-2004399,-2004376,-2004353,-2004331,-2004308,-2004285,-2004263,-2004240,-2004217,-2004194,-2004172,-2004149,-2004126,-2004103,-2004081,-2004058,-2004035,-2004012,-2003989,-2003967,-2003944,-2003921,-2003898,-2003875,-2003852,-2003829,-2003807,-2003784,-2003761,-2003738,-2003715,-2003692,-2003669,-2003646,-2003623,-2003600,-2003577,-2003554,-2003531,-2003508,-2003485,-2003462,-2003439,-2003416,-2003393,-2003370,-2003347,-2003324,-2003300,-2003277,-2003254,-2003231,-2003208,-2003185,-2003162,-2003139,-2003115,-2003092,-2003069,-2003046,-2003023,-2002999,-2002976,-2002953,-2002930,-2002906,-2002883,-2002860,-2002837,-2002813,-2002790,-2002767,-2002743,-2002720,-2002697,-2002673,-2002650,-2002627,-2002603,-2002580,-2002556,-2002533,-2002510,-2002486,-2002463,-2002439,-2002416,-2002392,-2002369,-2002345,-2002322,-2002298,-2002275,-2002251,-2002228,-2002204,-2002181,-2002157,-2002134,-2002110,-2002086,-2002063,-2002039,-2002016,-2001992,-2001968,-2001945,-2001921,-2001897,-2001874,-2001850,-2001826,-2001803,-2001779,-2001755,-2001732,-2001708,-2001684,-2001660,-2001637,-2001613,-2001589,-2001565,-2001541,-2001518,-2001494,-2001470,-2001446,-2001422,-2001398,-2001375,-2001351,-2001327,-2001303,-2001279,-2001255,-2001231,-2001207,-2001183,-2001159,-2001135,-2001111,-2001088,-2001064,-2001040,-2001016,-2000992,-2000968,-2000943,-2000919,-2000895,-2000871,-2000847,-2000823,-2000799,-2000775,-2000751,-2000727,-2000703,-2000679,-2000654,-2000630,-2000606,-2000582,-2000558,-2000534,-2000509,-2000485,-2000461,-2000437,-2000412,-2000388,-2000364,-2000340,-2000315,-2000291,-2000267,-2000243,-2000218,-2000194,-2000170,-2000145,-2000121,-2000097,-2000072,-2000048,-2000023,-1999999,-1999975,-1999950,-1999926,-1999901,-1999877,-1999852,-1999828,-1999804,-1999779,-1999755,-1999730,-1999706,-1999681,-1999657,-1999632,-1999607,-1999583,-1999558,-1999534,-1999509,-1999485,-1999460,-1999435,-1999411,-1999386,-1999362,-1999337,-1999312,-1999288,-1999263,-1999238,-1999214,-1999189,-1999164,-1999139,-1999115,-1999090,-1999065,-1999040,-1999016,-1998991,-1998966,-1998941,-1998917,-1998892,-1998867,-1998842,-1998817,-1998792,-1998768,-1998743,-1998718,-1998693,-1998668,-1998643,-1998618,-1998593,-1998568,-1998543,-1998518,-1998493,-1998469,-1998444,-1998419,-1998394,-1998369,-1998344,-1998319,-1998293,-1998268,-1998243,-1998218,-1998193,-1998168,-1998143,-1998118,-1998093,-1998068,-1998043,-1998017,-1997992,-1997967,-1997942,-1997917,-1997892,-1997866,-1997841,-1997816,-1997791,-1997766,-1997740,-1997715,-1997690,-1997665,-1997639,-1997614,-1997589,-1997563,-1997538,-1997513,-1997487,-1997462,-1997437,-1997411,-1997386,-1997361,-1997335,-1997310,-1997284,-1997259,-1997234,-1997208,-1997183,-1997157,-1997132,-1997106,-1997081,-1997055,-1997030,-1997004,-1996979,-1996953,-1996928,-1996902,-1996877,-1996851,-1996826,-1996800,-1996774,-1996749,-1996723,-1996698,-1996672,-1996646,-1996621,-1996595,-1996569,-1996544,-1996518,-1996492,-1996467,-1996441,-1996415,-1996389,-1996364,-1996338,-1996312,-1996286,-1996261,-1996235,-1996209,-1996183,-1996157,-1996132,-1996106,-1996080,-1996054,-1996028,-1996002,-1995977,-1995951,-1995925,-1995899,-1995873,-1995847,-1995821,-1995795,-1995769,-1995743,-1995717,-1995691,-1995665,-1995639,-1995613,-1995587,-1995561,-1995535,-1995509,-1995483,-1995457,-1995431,-1995405,-1995379,-1995353,-1995327,-1995300,-1995274,-1995248,-1995222,-1995196,-1995170,-1995143,-1995117,-1995091,-1995065,-1995039,-1995012,-1994986,-1994960,-1994934,-1994907,-1994881,-1994855,-1994829,-1994802,-1994776,-1994750,-1994723,-1994697,-1994671,-1994644,-1994618,-1994592,-1994565,-1994539,-1994512,-1994486,-1994460,-1994433,-1994407,-1994380,-1994354,-1994327,-1994301,-1994274,-1994248,-1994221,-1994195,-1994168,-1994142,-1994115,-1994089,-1994062,-1994036,-1994009,-1993983,-1993956,-1993929,-1993903,-1993876,-1993850,-1993823,-1993796,-1993770,-1993743,-1993716,-1993690,-1993663,-1993636,-1993609,-1993583,-1993556,-1993529,-1993502,-1993476,-1993449,-1993422,-1993395,-1993369,-1993342,-1993315,-1993288,-1993261,-1993234,-1993208,-1993181,-1993154,-1993127,-1993100,-1993073,-1993046,-1993019,-1992992,-1992966,-1992939,-1992912,-1992885,-1992858,-1992831,-1992804,-1992777,-1992750,-1992723,-1992696,-1992669,-1992642,-1992615,-1992587,-1992560,-1992533,-1992506,-1992479,-1992452,-1992425,-1992398,-1992371,-1992343,-1992316,-1992289,-1992262,-1992235,-1992208,-1992180,-1992153,-1992126,-1992099,-1992071,-1992044,-1992017,-1991990,-1991962,-1991935,-1991908,-1991880,-1991853,-1991826,-1991799,-1991771,-1991744,-1991716,-1991689,-1991662,-1991634,-1991607,-1991580,-1991552,-1991525,-1991497,-1991470,-1991442,-1991415,-1991387,-1991360,-1991332,-1991305,-1991277,-1991250,-1991222,-1991195,-1991167,-1991140,-1991112,-1991085,-1991057,-1991029,-1991002,-1990974,-1990947,-1990919,-1990891,-1990864,-1990836,-1990808,-1990781,-1990753,-1990725,-1990698,-1990670,-1990642,-1990614,-1990587,-1990559,-1990531,-1990503,-1990476,-1990448,-1990420,-1990392,-1990364,-1990337,-1990309,-1990281,-1990253,-1990225,-1990197,-1990169,-1990142,-1990114,-1990086,-1990058,-1990030,-1990002,-1989974,-1989946,-1989918,-1989890,-1989862,-1989834,-1989806,-1989778,-1989750,-1989722,-1989694,-1989666,-1989638,-1989610,-1989582,-1989554,-1989526,-1989498,-1989469,-1989441,-1989413,-1989385,-1989357,-1989329,-1989301,-1989272,-1989244,-1989216,-1989188,-1989160,-1989131,-1989103,-1989075,-1989047,-1989018,-1988990,-1988962,-1988934,-1988905,-1988877,-1988849,-1988820,-1988792,-1988764,-1988735,-1988707,-1988679,-1988650,-1988622,-1988593,-1988565,-1988537,-1988508,-1988480,-1988451,-1988423,-1988394,-1988366,-1988337,-1988309,-1988280,-1988252,-1988223,-1988195,-1988166,-1988138,-1988109,-1988081,-1988052,-1988023,-1987995,-1987966,-1987938,-1987909,-1987880,-1987852,-1987823,-1987795,-1987766,-1987737,-1987708,-1987680,-1987651,-1987622,-1987594,-1987565,-1987536,-1987507,-1987479,-1987450,-1987421,-1987392,-1987364,-1987335,-1987306,-1987277,-1987248,-1987219,-1987191,-1987162,-1987133,-1987104,-1987075,-1987046,-1987017,-1986988,-1986959,-1986931,-1986902,-1986873,-1986844,-1986815,-1986786,-1986757,-1986728,-1986699,-1986670,-1986641,-1986612,-1986583,-1986554,-1986524,-1986495,-1986466,-1986437,-1986408,-1986379,-1986350,-1986321,-1986292,-1986262,-1986233,-1986204,-1986175,-1986146,-1986117,-1986087,-1986058,-1986029,-1986000,-1985971,-1985941,-1985912,-1985883,-1985853,-1985824,-1985795,-1985766,-1985736,-1985707,-1985678,-1985648,-1985619,-1985590,-1985560,-1985531,-1985501,-1985472,-1985443,-1985413,-1985384,-1985354,-1985325,-1985295,-1985266,-1985237,-1985207,-1985178,-1985148,-1985119,-1985089,-1985060,-1985030,-1985000,-1984971,-1984941,-1984912,-1984882,-1984853,-1984823,-1984793,-1984764,-1984734,-1984705,-1984675,-1984645,-1984616,-1984586,-1984556,-1984527,-1984497,-1984467,-1984437,-1984408,-1984378,-1984348,-1984318,-1984289,-1984259,-1984229,-1984199,-1984170,-1984140,-1984110,-1984080,-1984050,-1984020,-1983991,-1983961,-1983931,-1983901,-1983871,-1983841,-1983811,-1983781,-1983751,-1983721,-1983691,-1983661,-1983632,-1983602,-1983572,-1983542,-1983512,-1983482,-1983452,-1983421,-1983391,-1983361,-1983331,-1983301,-1983271,-1983241,-1983211,-1983181,-1983151,-1983121,-1983091,-1983060,-1983030,-1983000,-1982970,-1982940,-1982910,-1982879,-1982849,-1982819,-1982789,-1982758,-1982728,-1982698,-1982668,-1982637,-1982607,-1982577,-1982547,-1982516,-1982486,-1982456,-1982425,-1982395,-1982365,-1982334,-1982304,-1982273,-1982243,-1982213,-1982182,-1982152,-1982121,-1982091,-1982061,-1982030,-1982000,-1981969,-1981939,-1981908,-1981878,-1981847,-1981817,-1981786,-1981756,-1981725,-1981694,-1981664,-1981633,-1981603,-1981572,-1981542,-1981511,-1981480,-1981450,-1981419,-1981388,-1981358,-1981327,-1981296,-1981266,-1981235,-1981204,-1981174,-1981143,-1981112,-1981081,-1981051,-1981020,-1980989,-1980958,-1980928,-1980897,-1980866,-1980835,-1980804,-1980773,-1980743,-1980712,-1980681,-1980650,-1980619,-1980588,-1980557,-1980526,-1980496,-1980465,-1980434,-1980403,-1980372,-1980341,-1980310,-1980279,-1980248,-1980217,-1980186,-1980155,-1980124,-1980093,-1980062,-1980031,-1980000,-1979969,-1979937,-1979906,-1979875,-1979844,-1979813,-1979782,-1979751,-1979720,-1979688,-1979657,-1979626,-1979595,-1979564,-1979533,-1979501,-1979470,-1979439,-1979408,-1979376,-1979345,-1979314,-1979283,-1979251,-1979220,-1979189,-1979157,-1979126,-1979095,-1979063,-1979032,-1979001,-1978969,-1978938,-1978907,-1978875,-1978844,-1978812,-1978781,-1978750,-1978718,-1978687,-1978655,-1978624,-1978592,-1978561,-1978529,-1978498,-1978466,-1978435,-1978403,-1978372,-1978340,-1978309,-1978277,-1978245,-1978214,-1978182,-1978151,-1978119,-1978087,-1978056,-1978024,-1977992,-1977961,-1977929,-1977897,-1977866,-1977834,-1977802,-1977771,-1977739,-1977707,-1977675,-1977644,-1977612,-1977580,-1977548,-1977517,-1977485,-1977453,-1977421,-1977389,-1977357,-1977326,-1977294,-1977262,-1977230,-1977198,-1977166,-1977134,-1977102,-1977071,-1977039,-1977007,-1976975,-1976943,-1976911,-1976879,-1976847,-1976815,-1976783,-1976751,-1976719,-1976687,-1976655,-1976623,-1976591,-1976559,-1976526,-1976494,-1976462,-1976430,-1976398,-1976366,-1976334,-1976302,-1976270,-1976237,-1976205,-1976173,-1976141,-1976109,-1976076,-1976044,-1976012,-1975980,-1975948,-1975915,-1975883,-1975851,-1975819,-1975786,-1975754,-1975722,-1975689,-1975657,-1975625,-1975592,-1975560,-1975528,-1975495,-1975463,-1975430,-1975398,-1975366,-1975333,-1975301,-1975268,-1975236,-1975204,-1975171,-1975139,-1975106,-1975074,-1975041,-1975009,-1974976,-1974944,-1974911,-1974878,-1974846,-1974813,-1974781,-1974748,-1974716,-1974683,-1974650,-1974618,-1974585,-1974553,-1974520,-1974487,-1974455,-1974422,-1974389,-1974357,-1974324,-1974291,-1974258,-1974226,-1974193,-1974160,-1974127,-1974095,-1974062,-1974029,-1973996,-1973964,-1973931,-1973898,-1973865,-1973832,-1973799,-1973767,-1973734,-1973701,-1973668,-1973635,-1973602,-1973569,-1973536,-1973503,-1973470,-1973438,-1973405,-1973372,-1973339,-1973306,-1973273,-1973240,-1973207,-1973174,-1973141,-1973108,-1973074,-1973041,-1973008,-1972975,-1972942,-1972909,-1972876,-1972843,-1972810,-1972777,-1972744,-1972710,-1972677,-1972644,-1972611,-1972578,-1972544,-1972511,-1972478,-1972445,-1972412,-1972378,-1972345,-1972312,-1972279,-1972245,-1972212,-1972179,-1972145,-1972112,-1972079,-1972045,-1972012,-1971979,-1971945,-1971912,-1971879,-1971845,-1971812,-1971778,-1971745,-1971712,-1971678,-1971645,-1971611,-1971578,-1971544,-1971511,-1971477,-1971444,-1971410,-1971377,-1971343,-1971310,-1971276,-1971243,-1971209,-1971176,-1971142,-1971108,-1971075,-1971041,-1971008,-1970974,-1970940,-1970907,-1970873,-1970839,-1970806,-1970772,-1970738,-1970705,-1970671,-1970637,-1970604,-1970570,-1970536,-1970502,-1970469,-1970435,-1970401,-1970367,-1970333,-1970300,-1970266,-1970232,-1970198,-1970164,-1970130,-1970097,-1970063,-1970029,-1969995,-1969961,-1969927,-1969893,-1969859,-1969825,-1969791,-1969757,-1969723,-1969689,-1969655,-1969621,-1969587,-1969553,-1969519,-1969485,-1969451,-1969417,-1969383,-1969349,-1969315,-1969281,-1969247,-1969213,-1969179,-1969145,-1969110,-1969076,-1969042,-1969008,-1968974,-1968940,-1968906,-1968871,-1968837,-1968803,-1968769,-1968734,-1968700,-1968666,-1968632,-1968597,-1968563,-1968529,-1968495,-1968460,-1968426,-1968392,-1968357,-1968323,-1968289,-1968254,-1968220,-1968186,-1968151,-1968117,-1968082,-1968048,-1968014,-1967979,-1967945,-1967910,-1967876,-1967841,-1967807,-1967772,-1967738,-1967703,-1967669,-1967634,-1967600,-1967565,-1967531,-1967496,-1967462,-1967427,-1967392,-1967358,-1967323,-1967289,-1967254,-1967219,-1967185,-1967150,-1967115,-1967081,-1967046,-1967011,-1966977,-1966942,-1966907,-1966872,-1966838,-1966803,-1966768,-1966733,-1966699,-1966664,-1966629,-1966594,-1966560,-1966525,-1966490,-1966455,-1966420,-1966385,-1966351,-1966316,-1966281,-1966246,-1966211,-1966176,-1966141,-1966106,-1966071,-1966036,-1966001,-1965966,-1965931,-1965897,-1965862,-1965827,-1965792,-1965756,-1965721,-1965686,-1965651,-1965616,-1965581,-1965546,-1965511,-1965476,-1965441,-1965406,-1965371,-1965336,-1965300,-1965265,-1965230,-1965195,-1965160,-1965125,-1965089,-1965054,-1965019,-1964984,-1964949,-1964913,-1964878,-1964843,-1964808,-1964772,-1964737,-1964702,-1964666,-1964631,-1964596,-1964561,-1964525,-1964490,-1964454,-1964419,-1964384,-1964348,-1964313,-1964278,-1964242,-1964207,-1964171,-1964136,-1964100,-1964065,-1964030,-1963994,-1963959,-1963923,-1963888,-1963852,-1963817,-1963781,-1963745,-1963710,-1963674,-1963639,-1963603,-1963568,-1963532,-1963496,-1963461,-1963425,-1963390,-1963354,-1963318,-1963283,-1963247,-1963211,-1963176,-1963140,-1963104,-1963069,-1963033,-1962997,-1962961,-1962926,-1962890,-1962854,-1962818,-1962783,-1962747,-1962711,-1962675,-1962639,-1962603,-1962568,-1962532,-1962496,-1962460,-1962424,-1962388,-1962352,-1962317,-1962281,-1962245,-1962209,-1962173,-1962137,-1962101,-1962065,-1962029,-1961993,-1961957,-1961921,-1961885,-1961849,-1961813,-1961777,-1961741,-1961705,-1961669,-1961633,-1961597,-1961560,-1961524,-1961488,-1961452,-1961416,-1961380,-1961344,-1961308,-1961271,-1961235,-1961199,-1961163,-1961127,-1961090,-1961054,-1961018,-1960982,-1960946,-1960909,-1960873,-1960837,-1960800,-1960764,-1960728,-1960692,-1960655,-1960619,-1960583,-1960546,-1960510,-1960473,-1960437,-1960401,-1960364,-1960328,-1960291,-1960255,-1960219,-1960182,-1960146,-1960109,-1960073,-1960036,-1960000,-1959963,-1959927,-1959890,-1959854,-1959817,-1959781,-1959744,-1959708,-1959671,-1959635,-1959598,-1959561,-1959525,-1959488,-1959451,-1959415,-1959378,-1959342,-1959305,-1959268,-1959232,-1959195,-1959158,-1959121,-1959085,-1959048,-1959011,-1958975,-1958938,-1958901,-1958864,-1958828,-1958791,-1958754,-1958717,-1958680,-1958644,-1958607,-1958570,-1958533,-1958496,-1958459,-1958422,-1958386,-1958349,-1958312,-1958275,-1958238,-1958201,-1958164,-1958127,-1958090,-1958053,-1958016,-1957979,-1957942,-1957905,-1957868,-1957831,-1957794,-1957757,-1957720,-1957683,-1957646,-1957609,-1957572,-1957535,-1957498,-1957460,-1957423,-1957386,-1957349,-1957312,-1957275,-1957238,-1957200,-1957163,-1957126,-1957089,-1957052,-1957014,-1956977,-1956940,-1956903,-1956865,-1956828,-1956791,-1956754,-1956716,-1956679,-1956642,-1956604,-1956567,-1956530,-1956492,-1956455,-1956418,-1956380,-1956343,-1956305,-1956268,-1956231,-1956193,-1956156,-1956118,-1956081,-1956043,-1956006,-1955968,-1955931,-1955893,-1955856,-1955818,-1955781,-1955743,-1955706,-1955668,-1955631,-1955593,-1955556,-1955518,-1955480,-1955443,-1955405,-1955368,-1955330,-1955292,-1955255,-1955217,-1955179,-1955142,-1955104,-1955066,-1955029,-1954991,-1954953,-1954915,-1954878,-1954840,-1954802,-1954764,-1954727,-1954689,-1954651,-1954613,-1954575,-1954538,-1954500,-1954462,-1954424,-1954386,-1954348,-1954310,-1954273,-1954235,-1954197,-1954159,-1954121,-1954083,-1954045,-1954007,-1953969,-1953931,-1953893,-1953855,-1953817,-1953779,-1953741,-1953703,-1953665,-1953627,-1953589,-1953551,-1953513,-1953475,-1953437,-1953399,-1953361,-1953322,-1953284,-1953246,-1953208,-1953170,-1953132,-1953094,-1953055,-1953017,-1952979,-1952941,-1952903,-1952864,-1952826,-1952788,-1952750,-1952711,-1952673,-1952635,-1952597,-1952558,-1952520,-1952482,-1952443,-1952405,-1952367,-1952328,-1952290,-1952252,-1952213,-1952175,-1952136,-1952098,-1952060,-1952021,-1951983,-1951944,-1951906,-1951867,-1951829,-1951790);
signal constA1 : signed(w_coef-1 downto 0):= to_signed(-2079063,w_coef);
signal bp1_out : signed(W_in-1 downto 0) := (others =>'0');
signal BP_out : signed(W_in-1 downto 0) := (others =>'0');
signal data_out_temp:  signed(W_in-1 downto 0) := (others =>'0');
signal BW_clk : std_logic := '0';
signal newCLK : std_logic := '0';
signal count_int : integer:= 8000 ;

signal WahWah_EN : std_logic := '0';
begin

process(clk_50,nReset)
begin
if(rising_edge(clk_50)) then
	IF filterid(7 DOWNTO 0) ="00010110"THEN --range value spi
		count_int <= to_integer(signed(fil_data));
	elsif filterid(7 downto 0) = "00010101"then -- on off range value
		if fil_data(0) =  '1' then
			WahWah_EN <= '1';
		elsif fil_data(0) = '0' then
			WahWah_EN <= '0';
		end if;
	END IF;
end if;
end process;


process(CLK_50,nReset) -- 4.91 Hz, 1000 count : 49.1 Hz
variable counter : integer := 0;
begin
if (nReset = '0') then
	counter := 0;
	newCLK <= '0';
elsif(rising_edge(CLK_50)) then
	counter := counter + 1;
	if (counter = count_int ) then 
		newCLK <= NOT newCLK;
		counter := 0;
	end if;
end if;
end process;


process(newCLK,nReset) 
variable counter : integer := 0;
variable direction: std_logic := '0';
begin
if (nReset = '0') then
	counter := 0;
	direction:= '0';
elsif (rising_edge(newCLK)) then
	if (direction = '0') then
		constA1 <= to_signed(A1(counter),w_coef);
		counter := counter + 1;
		if(counter = Arr_size) then
			direction := '1';
		end if;
	end if;
	if(direction = '1') then
		counter := counter -1;
		constA1 <= to_signed(A1(counter),w_coef);
		if(counter = 0) then
			direction := '0';
		end if;
	end if;
end if;
end process;

IIRDF_inst : IIRDF1_BW 
generic map(
   W_in => W_in,
	W_coef => W_coef,
	A0 => A0,
	A2 => A2,
	B0 => B0,
	B1 => B1,
	B2 => B2
)
port map(
	iCLK => CLK_50,          
	iRESET_N => nReset,      
	new_val => new_val,        
	IIR_in => data_in,                 
	IIR_out => bp1_out,         
   A1 => constA1
);

IIRDF2_inst : IIRDF1_BW 
generic map(
   W_in => W_in,
	W_coef => W_coef,
	A0 => A0,
	A2 => A2,
	B0 => B0,
	B1 => B1,
	B2 => B2
)
port map(
	iCLK => CLK_50,          
	iRESET_N => nReset,      
	new_val => new_val,        
	IIR_in => bp1_out,                 
	IIR_out => BP_out,         
   A1 => constA1
);

process(CLK_50,nReset)
begin
if nReset = '0' then
	data_out <= (others => '0');
elsif(rising_edge(CLK_50)) then
	if(new_val = '1') then
	if WahWah_EN = '0' then
		data_out <= data_in;
	elsif WahWah_EN = '1' then
		data_out <= resize((BP_out*4+data_in/2),data_out'length); -- previously BP_out*4 and data_in/2
	end if;
	end if;
end if;
end process;
end;