library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity WahWah_FX is
port (
	CLK_50		: in std_logic;
	nReset		: in std_logic;
	new_val		: in std_logic;       -- indicates a new input value, input from data_over
	data_in		: in signed (15 downto 0);         
	data_out		: out signed (15 downto 0);   -- Output
	WahWah_EN 	: in std_logic
);
end entity WahWah_FX;

architecture behaviour of WahWah_FX is
constant W_coef : integer := 20;
constant W_in : integer := 16;
constant Arr_size : integer := 20000;

component IIRDF1_BW is
generic (
    W_in : integer ;
	 W_coef : integer   
);
port (
	iCLK            : in std_logic;
	iRESET_N        : in std_logic;
	new_val         : in std_logic;       -- indicates a new input value, input from data_over
	IIR_in          : in signed (15 downto 0);   -- singed is expected             
	IIR_out         : out signed (15 downto 0);   -- Output

	B0 : in signed(W_coef-1 downto 0);  
   B1 : in signed(W_coef-1 downto 0);
   B2 : in signed(W_coef-1 downto 0);
   A0 : in signed(W_coef-1 downto 0);
   A1 : in signed(W_coef-1 downto 0);
   A2 : in signed(W_coef-1 downto 0)
);
end component;

type cA0_array_type is array (0 to Arr_size) of integer;  --626 length
signal A0 : cA0_array_type:=(others => 262144);

type cA1_array_type is array (0 to Arr_size) of integer;
signal A1 : cA1_array_type:=(-509990,-509989,-509989,-509988,-509987,-509987,-509986,-509986,-509985,-509985,-509984,-509984,-509983,-509983,-509982,-509981,-509981,-509980,-509980,-509979,-509979,-509978,-509978,-509977,-509977,-509976,-509975,-509975,-509974,-509974,-509973,-509973,-509972,-509972,-509971,-509970,-509970,-509969,-509969,-509968,-509968,-509967,-509967,-509966,-509965,-509965,-509964,-509964,-509963,-509963,-509962,-509962,-509961,-509960,-509960,-509959,-509959,-509958,-509958,-509957,-509957,-509956,-509956,-509955,-509954,-509954,-509953,-509953,-509952,-509952,-509951,-509950,-509950,-509949,-509949,-509948,-509948,-509947,-509947,-509946,-509945,-509945,-509944,-509944,-509943,-509943,-509942,-509942,-509941,-509940,-509940,-509939,-509939,-509938,-509938,-509937,-509937,-509936,-509935,-509935,-509934,-509934,-509933,-509933,-509932,-509931,-509931,-509930,-509930,-509929,-509929,-509928,-509928,-509927,-509926,-509926,-509925,-509925,-509924,-509924,-509923,-509922,-509922,-509921,-509921,-509920,-509920,-509919,-509919,-509918,-509917,-509917,-509916,-509916,-509915,-509915,-509914,-509913,-509913,-509912,-509912,-509911,-509911,-509910,-509909,-509909,-509908,-509908,-509907,-509907,-509906,-509906,-509905,-509904,-509904,-509903,-509903,-509902,-509902,-509901,-509900,-509900,-509899,-509899,-509898,-509898,-509897,-509896,-509896,-509895,-509895,-509894,-509894,-509893,-509892,-509892,-509891,-509891,-509890,-509890,-509889,-509888,-509888,-509887,-509887,-509886,-509886,-509885,-509884,-509884,-509883,-509883,-509882,-509882,-509881,-509880,-509880,-509879,-509879,-509878,-509878,-509877,-509876,-509876,-509875,-509875,-509874,-509874,-509873,-509872,-509872,-509871,-509871,-509870,-509869,-509869,-509868,-509868,-509867,-509867,-509866,-509865,-509865,-509864,-509864,-509863,-509863,-509862,-509861,-509861,-509860,-509860,-509859,-509859,-509858,-509857,-509857,-509856,-509856,-509855,-509854,-509854,-509853,-509853,-509852,-509852,-509851,-509850,-509850,-509849,-509849,-509848,-509847,-509847,-509846,-509846,-509845,-509845,-509844,-509843,-509843,-509842,-509842,-509841,-509840,-509840,-509839,-509839,-509838,-509838,-509837,-509836,-509836,-509835,-509835,-509834,-509833,-509833,-509832,-509832,-509831,-509831,-509830,-509829,-509829,-509828,-509828,-509827,-509826,-509826,-509825,-509825,-509824,-509824,-509823,-509822,-509822,-509821,-509821,-509820,-509819,-509819,-509818,-509818,-509817,-509816,-509816,-509815,-509815,-509814,-509814,-509813,-509812,-509812,-509811,-509811,-509810,-509809,-509809,-509808,-509808,-509807,-509806,-509806,-509805,-509805,-509804,-509803,-509803,-509802,-509802,-509801,-509801,-509800,-509799,-509799,-509798,-509798,-509797,-509796,-509796,-509795,-509795,-509794,-509793,-509793,-509792,-509792,-509791,-509790,-509790,-509789,-509789,-509788,-509787,-509787,-509786,-509786,-509785,-509784,-509784,-509783,-509783,-509782,-509782,-509781,-509780,-509780,-509779,-509779,-509778,-509777,-509777,-509776,-509776,-509775,-509774,-509774,-509773,-509773,-509772,-509771,-509771,-509770,-509770,-509769,-509768,-509768,-509767,-509767,-509766,-509765,-509765,-509764,-509764,-509763,-509762,-509762,-509761,-509761,-509760,-509759,-509759,-509758,-509758,-509757,-509756,-509756,-509755,-509755,-509754,-509753,-509753,-509752,-509751,-509751,-509750,-509750,-509749,-509748,-509748,-509747,-509747,-509746,-509745,-509745,-509744,-509744,-509743,-509742,-509742,-509741,-509741,-509740,-509739,-509739,-509738,-509738,-509737,-509736,-509736,-509735,-509735,-509734,-509733,-509733,-509732,-509732,-509731,-509730,-509730,-509729,-509728,-509728,-509727,-509727,-509726,-509725,-509725,-509724,-509724,-509723,-509722,-509722,-509721,-509721,-509720,-509719,-509719,-509718,-509717,-509717,-509716,-509716,-509715,-509714,-509714,-509713,-509713,-509712,-509711,-509711,-509710,-509710,-509709,-509708,-509708,-509707,-509706,-509706,-509705,-509705,-509704,-509703,-509703,-509702,-509702,-509701,-509700,-509700,-509699,-509698,-509698,-509697,-509697,-509696,-509695,-509695,-509694,-509694,-509693,-509692,-509692,-509691,-509690,-509690,-509689,-509689,-509688,-509687,-509687,-509686,-509686,-509685,-509684,-509684,-509683,-509682,-509682,-509681,-509681,-509680,-509679,-509679,-509678,-509677,-509677,-509676,-509676,-509675,-509674,-509674,-509673,-509672,-509672,-509671,-509671,-509670,-509669,-509669,-509668,-509668,-509667,-509666,-509666,-509665,-509664,-509664,-509663,-509663,-509662,-509661,-509661,-509660,-509659,-509659,-509658,-509658,-509657,-509656,-509656,-509655,-509654,-509654,-509653,-509653,-509652,-509651,-509651,-509650,-509649,-509649,-509648,-509648,-509647,-509646,-509646,-509645,-509644,-509644,-509643,-509643,-509642,-509641,-509641,-509640,-509639,-509639,-509638,-509637,-509637,-509636,-509636,-509635,-509634,-509634,-509633,-509632,-509632,-509631,-509631,-509630,-509629,-509629,-509628,-509627,-509627,-509626,-509626,-509625,-509624,-509624,-509623,-509622,-509622,-509621,-509620,-509620,-509619,-509619,-509618,-509617,-509617,-509616,-509615,-509615,-509614,-509614,-509613,-509612,-509612,-509611,-509610,-509610,-509609,-509608,-509608,-509607,-509607,-509606,-509605,-509605,-509604,-509603,-509603,-509602,-509601,-509601,-509600,-509600,-509599,-509598,-509598,-509597,-509596,-509596,-509595,-509594,-509594,-509593,-509593,-509592,-509591,-509591,-509590,-509589,-509589,-509588,-509587,-509587,-509586,-509585,-509585,-509584,-509584,-509583,-509582,-509582,-509581,-509580,-509580,-509579,-509578,-509578,-509577,-509576,-509576,-509575,-509575,-509574,-509573,-509573,-509572,-509571,-509571,-509570,-509569,-509569,-509568,-509567,-509567,-509566,-509566,-509565,-509564,-509564,-509563,-509562,-509562,-509561,-509560,-509560,-509559,-509558,-509558,-509557,-509557,-509556,-509555,-509555,-509554,-509553,-509553,-509552,-509551,-509551,-509550,-509549,-509549,-509548,-509547,-509547,-509546,-509546,-509545,-509544,-509544,-509543,-509542,-509542,-509541,-509540,-509540,-509539,-509538,-509538,-509537,-509536,-509536,-509535,-509534,-509534,-509533,-509533,-509532,-509531,-509531,-509530,-509529,-509529,-509528,-509527,-509527,-509526,-509525,-509525,-509524,-509523,-509523,-509522,-509521,-509521,-509520,-509519,-509519,-509518,-509518,-509517,-509516,-509516,-509515,-509514,-509514,-509513,-509512,-509512,-509511,-509510,-509510,-509509,-509508,-509508,-509507,-509506,-509506,-509505,-509504,-509504,-509503,-509502,-509502,-509501,-509500,-509500,-509499,-509498,-509498,-509497,-509497,-509496,-509495,-509495,-509494,-509493,-509493,-509492,-509491,-509491,-509490,-509489,-509489,-509488,-509487,-509487,-509486,-509485,-509485,-509484,-509483,-509483,-509482,-509481,-509481,-509480,-509479,-509479,-509478,-509477,-509477,-509476,-509475,-509475,-509474,-509473,-509473,-509472,-509471,-509471,-509470,-509469,-509469,-509468,-509467,-509467,-509466,-509465,-509465,-509464,-509463,-509463,-509462,-509461,-509461,-509460,-509459,-509459,-509458,-509457,-509457,-509456,-509455,-509455,-509454,-509453,-509453,-509452,-509451,-509451,-509450,-509449,-509449,-509448,-509447,-509447,-509446,-509445,-509445,-509444,-509443,-509443,-509442,-509441,-509441,-509440,-509439,-509439,-509438,-509437,-509437,-509436,-509435,-509435,-509434,-509433,-509433,-509432,-509431,-509431,-509430,-509429,-509429,-509428,-509427,-509427,-509426,-509425,-509425,-509424,-509423,-509423,-509422,-509421,-509421,-509420,-509419,-509419,-509418,-509417,-509416,-509416,-509415,-509414,-509414,-509413,-509412,-509412,-509411,-509410,-509410,-509409,-509408,-509408,-509407,-509406,-509406,-509405,-509404,-509404,-509403,-509402,-509402,-509401,-509400,-509400,-509399,-509398,-509398,-509397,-509396,-509395,-509395,-509394,-509393,-509393,-509392,-509391,-509391,-509390,-509389,-509389,-509388,-509387,-509387,-509386,-509385,-509385,-509384,-509383,-509383,-509382,-509381,-509381,-509380,-509379,-509378,-509378,-509377,-509376,-509376,-509375,-509374,-509374,-509373,-509372,-509372,-509371,-509370,-509370,-509369,-509368,-509368,-509367,-509366,-509365,-509365,-509364,-509363,-509363,-509362,-509361,-509361,-509360,-509359,-509359,-509358,-509357,-509357,-509356,-509355,-509354,-509354,-509353,-509352,-509352,-509351,-509350,-509350,-509349,-509348,-509348,-509347,-509346,-509346,-509345,-509344,-509343,-509343,-509342,-509341,-509341,-509340,-509339,-509339,-509338,-509337,-509337,-509336,-509335,-509334,-509334,-509333,-509332,-509332,-509331,-509330,-509330,-509329,-509328,-509328,-509327,-509326,-509325,-509325,-509324,-509323,-509323,-509322,-509321,-509321,-509320,-509319,-509319,-509318,-509317,-509316,-509316,-509315,-509314,-509314,-509313,-509312,-509312,-509311,-509310,-509310,-509309,-509308,-509307,-509307,-509306,-509305,-509305,-509304,-509303,-509303,-509302,-509301,-509300,-509300,-509299,-509298,-509298,-509297,-509296,-509296,-509295,-509294,-509293,-509293,-509292,-509291,-509291,-509290,-509289,-509289,-509288,-509287,-509286,-509286,-509285,-509284,-509284,-509283,-509282,-509282,-509281,-509280,-509279,-509279,-509278,-509277,-509277,-509276,-509275,-509275,-509274,-509273,-509272,-509272,-509271,-509270,-509270,-509269,-509268,-509267,-509267,-509266,-509265,-509265,-509264,-509263,-509263,-509262,-509261,-509260,-509260,-509259,-509258,-509258,-509257,-509256,-509255,-509255,-509254,-509253,-509253,-509252,-509251,-509251,-509250,-509249,-509248,-509248,-509247,-509246,-509246,-509245,-509244,-509243,-509243,-509242,-509241,-509241,-509240,-509239,-509238,-509238,-509237,-509236,-509236,-509235,-509234,-509234,-509233,-509232,-509231,-509231,-509230,-509229,-509229,-509228,-509227,-509226,-509226,-509225,-509224,-509224,-509223,-509222,-509221,-509221,-509220,-509219,-509219,-509218,-509217,-509216,-509216,-509215,-509214,-509214,-509213,-509212,-509211,-509211,-509210,-509209,-509209,-509208,-509207,-509206,-509206,-509205,-509204,-509204,-509203,-509202,-509201,-509201,-509200,-509199,-509199,-509198,-509197,-509196,-509196,-509195,-509194,-509193,-509193,-509192,-509191,-509191,-509190,-509189,-509188,-509188,-509187,-509186,-509186,-509185,-509184,-509183,-509183,-509182,-509181,-509181,-509180,-509179,-509178,-509178,-509177,-509176,-509175,-509175,-509174,-509173,-509173,-509172,-509171,-509170,-509170,-509169,-509168,-509168,-509167,-509166,-509165,-509165,-509164,-509163,-509162,-509162,-509161,-509160,-509160,-509159,-509158,-509157,-509157,-509156,-509155,-509154,-509154,-509153,-509152,-509152,-509151,-509150,-509149,-509149,-509148,-509147,-509146,-509146,-509145,-509144,-509144,-509143,-509142,-509141,-509141,-509140,-509139,-509138,-509138,-509137,-509136,-509136,-509135,-509134,-509133,-509133,-509132,-509131,-509130,-509130,-509129,-509128,-509128,-509127,-509126,-509125,-509125,-509124,-509123,-509122,-509122,-509121,-509120,-509119,-509119,-509118,-509117,-509117,-509116,-509115,-509114,-509114,-509113,-509112,-509111,-509111,-509110,-509109,-509108,-509108,-509107,-509106,-509106,-509105,-509104,-509103,-509103,-509102,-509101,-509100,-509100,-509099,-509098,-509097,-509097,-509096,-509095,-509094,-509094,-509093,-509092,-509092,-509091,-509090,-509089,-509089,-509088,-509087,-509086,-509086,-509085,-509084,-509083,-509083,-509082,-509081,-509080,-509080,-509079,-509078,-509077,-509077,-509076,-509075,-509075,-509074,-509073,-509072,-509072,-509071,-509070,-509069,-509069,-509068,-509067,-509066,-509066,-509065,-509064,-509063,-509063,-509062,-509061,-509060,-509060,-509059,-509058,-509057,-509057,-509056,-509055,-509054,-509054,-509053,-509052,-509051,-509051,-509050,-509049,-509048,-509048,-509047,-509046,-509046,-509045,-509044,-509043,-509043,-509042,-509041,-509040,-509040,-509039,-509038,-509037,-509037,-509036,-509035,-509034,-509034,-509033,-509032,-509031,-509031,-509030,-509029,-509028,-509028,-509027,-509026,-509025,-509025,-509024,-509023,-509022,-509022,-509021,-509020,-509019,-509019,-509018,-509017,-509016,-509016,-509015,-509014,-509013,-509013,-509012,-509011,-509010,-509010,-509009,-509008,-509007,-509007,-509006,-509005,-509004,-509004,-509003,-509002,-509001,-509000,-509000,-508999,-508998,-508997,-508997,-508996,-508995,-508994,-508994,-508993,-508992,-508991,-508991,-508990,-508989,-508988,-508988,-508987,-508986,-508985,-508985,-508984,-508983,-508982,-508982,-508981,-508980,-508979,-508979,-508978,-508977,-508976,-508976,-508975,-508974,-508973,-508972,-508972,-508971,-508970,-508969,-508969,-508968,-508967,-508966,-508966,-508965,-508964,-508963,-508963,-508962,-508961,-508960,-508960,-508959,-508958,-508957,-508957,-508956,-508955,-508954,-508953,-508953,-508952,-508951,-508950,-508950,-508949,-508948,-508947,-508947,-508946,-508945,-508944,-508944,-508943,-508942,-508941,-508940,-508940,-508939,-508938,-508937,-508937,-508936,-508935,-508934,-508934,-508933,-508932,-508931,-508931,-508930,-508929,-508928,-508927,-508927,-508926,-508925,-508924,-508924,-508923,-508922,-508921,-508921,-508920,-508919,-508918,-508917,-508917,-508916,-508915,-508914,-508914,-508913,-508912,-508911,-508911,-508910,-508909,-508908,-508907,-508907,-508906,-508905,-508904,-508904,-508903,-508902,-508901,-508900,-508900,-508899,-508898,-508897,-508897,-508896,-508895,-508894,-508894,-508893,-508892,-508891,-508890,-508890,-508889,-508888,-508887,-508887,-508886,-508885,-508884,-508883,-508883,-508882,-508881,-508880,-508880,-508879,-508878,-508877,-508876,-508876,-508875,-508874,-508873,-508873,-508872,-508871,-508870,-508869,-508869,-508868,-508867,-508866,-508866,-508865,-508864,-508863,-508862,-508862,-508861,-508860,-508859,-508859,-508858,-508857,-508856,-508855,-508855,-508854,-508853,-508852,-508852,-508851,-508850,-508849,-508848,-508848,-508847,-508846,-508845,-508845,-508844,-508843,-508842,-508841,-508841,-508840,-508839,-508838,-508837,-508837,-508836,-508835,-508834,-508834,-508833,-508832,-508831,-508830,-508830,-508829,-508828,-508827,-508827,-508826,-508825,-508824,-508823,-508823,-508822,-508821,-508820,-508819,-508819,-508818,-508817,-508816,-508816,-508815,-508814,-508813,-508812,-508812,-508811,-508810,-508809,-508808,-508808,-508807,-508806,-508805,-508804,-508804,-508803,-508802,-508801,-508801,-508800,-508799,-508798,-508797,-508797,-508796,-508795,-508794,-508793,-508793,-508792,-508791,-508790,-508789,-508789,-508788,-508787,-508786,-508785,-508785,-508784,-508783,-508782,-508782,-508781,-508780,-508779,-508778,-508778,-508777,-508776,-508775,-508774,-508774,-508773,-508772,-508771,-508770,-508770,-508769,-508768,-508767,-508766,-508766,-508765,-508764,-508763,-508762,-508762,-508761,-508760,-508759,-508758,-508758,-508757,-508756,-508755,-508754,-508754,-508753,-508752,-508751,-508751,-508750,-508749,-508748,-508747,-508747,-508746,-508745,-508744,-508743,-508743,-508742,-508741,-508740,-508739,-508739,-508738,-508737,-508736,-508735,-508735,-508734,-508733,-508732,-508731,-508731,-508730,-508729,-508728,-508727,-508726,-508726,-508725,-508724,-508723,-508722,-508722,-508721,-508720,-508719,-508718,-508718,-508717,-508716,-508715,-508714,-508714,-508713,-508712,-508711,-508710,-508710,-508709,-508708,-508707,-508706,-508706,-508705,-508704,-508703,-508702,-508702,-508701,-508700,-508699,-508698,-508698,-508697,-508696,-508695,-508694,-508693,-508693,-508692,-508691,-508690,-508689,-508689,-508688,-508687,-508686,-508685,-508685,-508684,-508683,-508682,-508681,-508681,-508680,-508679,-508678,-508677,-508676,-508676,-508675,-508674,-508673,-508672,-508672,-508671,-508670,-508669,-508668,-508668,-508667,-508666,-508665,-508664,-508663,-508663,-508662,-508661,-508660,-508659,-508659,-508658,-508657,-508656,-508655,-508655,-508654,-508653,-508652,-508651,-508650,-508650,-508649,-508648,-508647,-508646,-508646,-508645,-508644,-508643,-508642,-508641,-508641,-508640,-508639,-508638,-508637,-508637,-508636,-508635,-508634,-508633,-508632,-508632,-508631,-508630,-508629,-508628,-508628,-508627,-508626,-508625,-508624,-508623,-508623,-508622,-508621,-508620,-508619,-508619,-508618,-508617,-508616,-508615,-508614,-508614,-508613,-508612,-508611,-508610,-508610,-508609,-508608,-508607,-508606,-508605,-508605,-508604,-508603,-508602,-508601,-508600,-508600,-508599,-508598,-508597,-508596,-508596,-508595,-508594,-508593,-508592,-508591,-508591,-508590,-508589,-508588,-508587,-508586,-508586,-508585,-508584,-508583,-508582,-508582,-508581,-508580,-508579,-508578,-508577,-508577,-508576,-508575,-508574,-508573,-508572,-508572,-508571,-508570,-508569,-508568,-508567,-508567,-508566,-508565,-508564,-508563,-508562,-508562,-508561,-508560,-508559,-508558,-508557,-508557,-508556,-508555,-508554,-508553,-508552,-508552,-508551,-508550,-508549,-508548,-508548,-508547,-508546,-508545,-508544,-508543,-508543,-508542,-508541,-508540,-508539,-508538,-508538,-508537,-508536,-508535,-508534,-508533,-508533,-508532,-508531,-508530,-508529,-508528,-508527,-508527,-508526,-508525,-508524,-508523,-508522,-508522,-508521,-508520,-508519,-508518,-508517,-508517,-508516,-508515,-508514,-508513,-508512,-508512,-508511,-508510,-508509,-508508,-508507,-508507,-508506,-508505,-508504,-508503,-508502,-508502,-508501,-508500,-508499,-508498,-508497,-508496,-508496,-508495,-508494,-508493,-508492,-508491,-508491,-508490,-508489,-508488,-508487,-508486,-508486,-508485,-508484,-508483,-508482,-508481,-508480,-508480,-508479,-508478,-508477,-508476,-508475,-508475,-508474,-508473,-508472,-508471,-508470,-508470,-508469,-508468,-508467,-508466,-508465,-508464,-508464,-508463,-508462,-508461,-508460,-508459,-508459,-508458,-508457,-508456,-508455,-508454,-508453,-508453,-508452,-508451,-508450,-508449,-508448,-508448,-508447,-508446,-508445,-508444,-508443,-508442,-508442,-508441,-508440,-508439,-508438,-508437,-508436,-508436,-508435,-508434,-508433,-508432,-508431,-508431,-508430,-508429,-508428,-508427,-508426,-508425,-508425,-508424,-508423,-508422,-508421,-508420,-508419,-508419,-508418,-508417,-508416,-508415,-508414,-508413,-508413,-508412,-508411,-508410,-508409,-508408,-508407,-508407,-508406,-508405,-508404,-508403,-508402,-508401,-508401,-508400,-508399,-508398,-508397,-508396,-508396,-508395,-508394,-508393,-508392,-508391,-508390,-508390,-508389,-508388,-508387,-508386,-508385,-508384,-508383,-508383,-508382,-508381,-508380,-508379,-508378,-508377,-508377,-508376,-508375,-508374,-508373,-508372,-508371,-508371,-508370,-508369,-508368,-508367,-508366,-508365,-508365,-508364,-508363,-508362,-508361,-508360,-508359,-508359,-508358,-508357,-508356,-508355,-508354,-508353,-508352,-508352,-508351,-508350,-508349,-508348,-508347,-508346,-508346,-508345,-508344,-508343,-508342,-508341,-508340,-508340,-508339,-508338,-508337,-508336,-508335,-508334,-508333,-508333,-508332,-508331,-508330,-508329,-508328,-508327,-508327,-508326,-508325,-508324,-508323,-508322,-508321,-508320,-508320,-508319,-508318,-508317,-508316,-508315,-508314,-508314,-508313,-508312,-508311,-508310,-508309,-508308,-508307,-508307,-508306,-508305,-508304,-508303,-508302,-508301,-508300,-508300,-508299,-508298,-508297,-508296,-508295,-508294,-508293,-508293,-508292,-508291,-508290,-508289,-508288,-508287,-508286,-508286,-508285,-508284,-508283,-508282,-508281,-508280,-508279,-508279,-508278,-508277,-508276,-508275,-508274,-508273,-508272,-508272,-508271,-508270,-508269,-508268,-508267,-508266,-508265,-508265,-508264,-508263,-508262,-508261,-508260,-508259,-508258,-508258,-508257,-508256,-508255,-508254,-508253,-508252,-508251,-508251,-508250,-508249,-508248,-508247,-508246,-508245,-508244,-508243,-508243,-508242,-508241,-508240,-508239,-508238,-508237,-508236,-508236,-508235,-508234,-508233,-508232,-508231,-508230,-508229,-508229,-508228,-508227,-508226,-508225,-508224,-508223,-508222,-508221,-508221,-508220,-508219,-508218,-508217,-508216,-508215,-508214,-508213,-508213,-508212,-508211,-508210,-508209,-508208,-508207,-508206,-508206,-508205,-508204,-508203,-508202,-508201,-508200,-508199,-508198,-508198,-508197,-508196,-508195,-508194,-508193,-508192,-508191,-508190,-508190,-508189,-508188,-508187,-508186,-508185,-508184,-508183,-508182,-508182,-508181,-508180,-508179,-508178,-508177,-508176,-508175,-508174,-508174,-508173,-508172,-508171,-508170,-508169,-508168,-508167,-508166,-508165,-508165,-508164,-508163,-508162,-508161,-508160,-508159,-508158,-508157,-508157,-508156,-508155,-508154,-508153,-508152,-508151,-508150,-508149,-508148,-508148,-508147,-508146,-508145,-508144,-508143,-508142,-508141,-508140,-508140,-508139,-508138,-508137,-508136,-508135,-508134,-508133,-508132,-508131,-508131,-508130,-508129,-508128,-508127,-508126,-508125,-508124,-508123,-508122,-508122,-508121,-508120,-508119,-508118,-508117,-508116,-508115,-508114,-508113,-508113,-508112,-508111,-508110,-508109,-508108,-508107,-508106,-508105,-508104,-508104,-508103,-508102,-508101,-508100,-508099,-508098,-508097,-508096,-508095,-508095,-508094,-508093,-508092,-508091,-508090,-508089,-508088,-508087,-508086,-508086,-508085,-508084,-508083,-508082,-508081,-508080,-508079,-508078,-508077,-508076,-508076,-508075,-508074,-508073,-508072,-508071,-508070,-508069,-508068,-508067,-508066,-508066,-508065,-508064,-508063,-508062,-508061,-508060,-508059,-508058,-508057,-508056,-508056,-508055,-508054,-508053,-508052,-508051,-508050,-508049,-508048,-508047,-508046,-508046,-508045,-508044,-508043,-508042,-508041,-508040,-508039,-508038,-508037,-508036,-508036,-508035,-508034,-508033,-508032,-508031,-508030,-508029,-508028,-508027,-508026,-508026,-508025,-508024,-508023,-508022,-508021,-508020,-508019,-508018,-508017,-508016,-508015,-508015,-508014,-508013,-508012,-508011,-508010,-508009,-508008,-508007,-508006,-508005,-508004,-508004,-508003,-508002,-508001,-508000,-507999,-507998,-507997,-507996,-507995,-507994,-507993,-507993,-507992,-507991,-507990,-507989,-507988,-507987,-507986,-507985,-507984,-507983,-507982,-507982,-507981,-507980,-507979,-507978,-507977,-507976,-507975,-507974,-507973,-507972,-507971,-507970,-507970,-507969,-507968,-507967,-507966,-507965,-507964,-507963,-507962,-507961,-507960,-507959,-507958,-507958,-507957,-507956,-507955,-507954,-507953,-507952,-507951,-507950,-507949,-507948,-507947,-507946,-507946,-507945,-507944,-507943,-507942,-507941,-507940,-507939,-507938,-507937,-507936,-507935,-507934,-507933,-507933,-507932,-507931,-507930,-507929,-507928,-507927,-507926,-507925,-507924,-507923,-507922,-507921,-507920,-507920,-507919,-507918,-507917,-507916,-507915,-507914,-507913,-507912,-507911,-507910,-507909,-507908,-507907,-507907,-507906,-507905,-507904,-507903,-507902,-507901,-507900,-507899,-507898,-507897,-507896,-507895,-507894,-507893,-507893,-507892,-507891,-507890,-507889,-507888,-507887,-507886,-507885,-507884,-507883,-507882,-507881,-507880,-507879,-507879,-507878,-507877,-507876,-507875,-507874,-507873,-507872,-507871,-507870,-507869,-507868,-507867,-507866,-507865,-507864,-507864,-507863,-507862,-507861,-507860,-507859,-507858,-507857,-507856,-507855,-507854,-507853,-507852,-507851,-507850,-507849,-507849,-507848,-507847,-507846,-507845,-507844,-507843,-507842,-507841,-507840,-507839,-507838,-507837,-507836,-507835,-507834,-507833,-507833,-507832,-507831,-507830,-507829,-507828,-507827,-507826,-507825,-507824,-507823,-507822,-507821,-507820,-507819,-507818,-507817,-507817,-507816,-507815,-507814,-507813,-507812,-507811,-507810,-507809,-507808,-507807,-507806,-507805,-507804,-507803,-507802,-507801,-507800,-507799,-507799,-507798,-507797,-507796,-507795,-507794,-507793,-507792,-507791,-507790,-507789,-507788,-507787,-507786,-507785,-507784,-507783,-507782,-507781,-507781,-507780,-507779,-507778,-507777,-507776,-507775,-507774,-507773,-507772,-507771,-507770,-507769,-507768,-507767,-507766,-507765,-507764,-507763,-507762,-507762,-507761,-507760,-507759,-507758,-507757,-507756,-507755,-507754,-507753,-507752,-507751,-507750,-507749,-507748,-507747,-507746,-507745,-507744,-507743,-507742,-507741,-507741,-507740,-507739,-507738,-507737,-507736,-507735,-507734,-507733,-507732,-507731,-507730,-507729,-507728,-507727,-507726,-507725,-507724,-507723,-507722,-507721,-507720,-507719,-507719,-507718,-507717,-507716,-507715,-507714,-507713,-507712,-507711,-507710,-507709,-507708,-507707,-507706,-507705,-507704,-507703,-507702,-507701,-507700,-507699,-507698,-507697,-507696,-507696,-507695,-507694,-507693,-507692,-507691,-507690,-507689,-507688,-507687,-507686,-507685,-507684,-507683,-507682,-507681,-507680,-507679,-507678,-507677,-507676,-507675,-507674,-507673,-507672,-507671,-507670,-507669,-507669,-507668,-507667,-507666,-507665,-507664,-507663,-507662,-507661,-507660,-507659,-507658,-507657,-507656,-507655,-507654,-507653,-507652,-507651,-507650,-507649,-507648,-507647,-507646,-507645,-507644,-507643,-507642,-507641,-507640,-507640,-507639,-507638,-507637,-507636,-507635,-507634,-507633,-507632,-507631,-507630,-507629,-507628,-507627,-507626,-507625,-507624,-507623,-507622,-507621,-507620,-507619,-507618,-507617,-507616,-507615,-507614,-507613,-507612,-507611,-507610,-507609,-507608,-507607,-507606,-507606,-507605,-507604,-507603,-507602,-507601,-507600,-507599,-507598,-507597,-507596,-507595,-507594,-507593,-507592,-507591,-507590,-507589,-507588,-507587,-507586,-507585,-507584,-507583,-507582,-507581,-507580,-507579,-507578,-507577,-507576,-507575,-507574,-507573,-507572,-507571,-507570,-507569,-507568,-507567,-507566,-507565,-507564,-507563,-507563,-507562,-507561,-507560,-507559,-507558,-507557,-507556,-507555,-507554,-507553,-507552,-507551,-507550,-507549,-507548,-507547,-507546,-507545,-507544,-507543,-507542,-507541,-507540,-507539,-507538,-507537,-507536,-507535,-507534,-507533,-507532,-507531,-507530,-507529,-507528,-507527,-507526,-507525,-507524,-507523,-507522,-507521,-507520,-507519,-507518,-507517,-507516,-507515,-507514,-507513,-507512,-507511,-507510,-507509,-507508,-507507,-507506,-507505,-507504,-507503,-507502,-507501,-507500,-507500,-507499,-507498,-507497,-507496,-507495,-507494,-507493,-507492,-507491,-507490,-507489,-507488,-507487,-507486,-507485,-507484,-507483,-507482,-507481,-507480,-507479,-507478,-507477,-507476,-507475,-507474,-507473,-507472,-507471,-507470,-507469,-507468,-507467,-507466,-507465,-507464,-507463,-507462,-507461,-507460,-507459,-507458,-507457,-507456,-507455,-507454,-507453,-507452,-507451,-507450,-507449,-507448,-507447,-507446,-507445,-507444,-507443,-507442,-507441,-507440,-507439,-507438,-507437,-507436,-507435,-507434,-507433,-507432,-507431,-507430,-507429,-507428,-507427,-507426,-507425,-507424,-507423,-507422,-507421,-507420,-507419,-507418,-507417,-507416,-507415,-507414,-507413,-507412,-507411,-507410,-507409,-507408,-507407,-507406,-507405,-507404,-507403,-507402,-507401,-507400,-507399,-507398,-507397,-507396,-507395,-507394,-507393,-507392,-507391,-507390,-507389,-507388,-507387,-507386,-507385,-507384,-507383,-507382,-507381,-507380,-507379,-507378,-507377,-507376,-507375,-507374,-507373,-507372,-507371,-507370,-507369,-507368,-507367,-507366,-507365,-507364,-507363,-507362,-507361,-507360,-507359,-507358,-507357,-507356,-507355,-507354,-507353,-507352,-507351,-507350,-507349,-507348,-507347,-507346,-507345,-507344,-507343,-507342,-507341,-507340,-507339,-507338,-507337,-507336,-507335,-507334,-507332,-507331,-507330,-507329,-507328,-507327,-507326,-507325,-507324,-507323,-507322,-507321,-507320,-507319,-507318,-507317,-507316,-507315,-507314,-507313,-507312,-507311,-507310,-507309,-507308,-507307,-507306,-507305,-507304,-507303,-507302,-507301,-507300,-507299,-507298,-507297,-507296,-507295,-507294,-507293,-507292,-507291,-507290,-507289,-507288,-507287,-507286,-507285,-507284,-507283,-507282,-507281,-507280,-507279,-507278,-507277,-507276,-507275,-507274,-507273,-507272,-507271,-507270,-507268,-507267,-507266,-507265,-507264,-507263,-507262,-507261,-507260,-507259,-507258,-507257,-507256,-507255,-507254,-507253,-507252,-507251,-507250,-507249,-507248,-507247,-507246,-507245,-507244,-507243,-507242,-507241,-507240,-507239,-507238,-507237,-507236,-507235,-507234,-507233,-507232,-507231,-507230,-507229,-507228,-507227,-507226,-507225,-507223,-507222,-507221,-507220,-507219,-507218,-507217,-507216,-507215,-507214,-507213,-507212,-507211,-507210,-507209,-507208,-507207,-507206,-507205,-507204,-507203,-507202,-507201,-507200,-507199,-507198,-507197,-507196,-507195,-507194,-507193,-507192,-507191,-507190,-507189,-507187,-507186,-507185,-507184,-507183,-507182,-507181,-507180,-507179,-507178,-507177,-507176,-507175,-507174,-507173,-507172,-507171,-507170,-507169,-507168,-507167,-507166,-507165,-507164,-507163,-507162,-507161,-507160,-507159,-507158,-507157,-507155,-507154,-507153,-507152,-507151,-507150,-507149,-507148,-507147,-507146,-507145,-507144,-507143,-507142,-507141,-507140,-507139,-507138,-507137,-507136,-507135,-507134,-507133,-507132,-507131,-507130,-507129,-507127,-507126,-507125,-507124,-507123,-507122,-507121,-507120,-507119,-507118,-507117,-507116,-507115,-507114,-507113,-507112,-507111,-507110,-507109,-507108,-507107,-507106,-507105,-507104,-507103,-507101,-507100,-507099,-507098,-507097,-507096,-507095,-507094,-507093,-507092,-507091,-507090,-507089,-507088,-507087,-507086,-507085,-507084,-507083,-507082,-507081,-507080,-507079,-507077,-507076,-507075,-507074,-507073,-507072,-507071,-507070,-507069,-507068,-507067,-507066,-507065,-507064,-507063,-507062,-507061,-507060,-507059,-507058,-507057,-507055,-507054,-507053,-507052,-507051,-507050,-507049,-507048,-507047,-507046,-507045,-507044,-507043,-507042,-507041,-507040,-507039,-507038,-507037,-507036,-507035,-507033,-507032,-507031,-507030,-507029,-507028,-507027,-507026,-507025,-507024,-507023,-507022,-507021,-507020,-507019,-507018,-507017,-507016,-507015,-507013,-507012,-507011,-507010,-507009,-507008,-507007,-507006,-507005,-507004,-507003,-507002,-507001,-507000,-506999,-506998,-506997,-506996,-506994,-506993,-506992,-506991,-506990,-506989,-506988,-506987,-506986,-506985,-506984,-506983,-506982,-506981,-506980,-506979,-506978,-506977,-506975,-506974,-506973,-506972,-506971,-506970,-506969,-506968,-506967,-506966,-506965,-506964,-506963,-506962,-506961,-506960,-506959,-506957,-506956,-506955,-506954,-506953,-506952,-506951,-506950,-506949,-506948,-506947,-506946,-506945,-506944,-506943,-506942,-506940,-506939,-506938,-506937,-506936,-506935,-506934,-506933,-506932,-506931,-506930,-506929,-506928,-506927,-506926,-506925,-506923,-506922,-506921,-506920,-506919,-506918,-506917,-506916,-506915,-506914,-506913,-506912,-506911,-506910,-506909,-506907,-506906,-506905,-506904,-506903,-506902,-506901,-506900,-506899,-506898,-506897,-506896,-506895,-506894,-506892,-506891,-506890,-506889,-506888,-506887,-506886,-506885,-506884,-506883,-506882,-506881,-506880,-506879,-506878,-506876,-506875,-506874,-506873,-506872,-506871,-506870,-506869,-506868,-506867,-506866,-506865,-506864,-506863,-506861,-506860,-506859,-506858,-506857,-506856,-506855,-506854,-506853,-506852,-506851,-506850,-506849,-506847,-506846,-506845,-506844,-506843,-506842,-506841,-506840,-506839,-506838,-506837,-506836,-506835,-506834,-506832,-506831,-506830,-506829,-506828,-506827,-506826,-506825,-506824,-506823,-506822,-506821,-506820,-506818,-506817,-506816,-506815,-506814,-506813,-506812,-506811,-506810,-506809,-506808,-506807,-506805,-506804,-506803,-506802,-506801,-506800,-506799,-506798,-506797,-506796,-506795,-506794,-506793,-506791,-506790,-506789,-506788,-506787,-506786,-506785,-506784,-506783,-506782,-506781,-506780,-506778,-506777,-506776,-506775,-506774,-506773,-506772,-506771,-506770,-506769,-506768,-506767,-506765,-506764,-506763,-506762,-506761,-506760,-506759,-506758,-506757,-506756,-506755,-506753,-506752,-506751,-506750,-506749,-506748,-506747,-506746,-506745,-506744,-506743,-506742,-506740,-506739,-506738,-506737,-506736,-506735,-506734,-506733,-506732,-506731,-506730,-506728,-506727,-506726,-506725,-506724,-506723,-506722,-506721,-506720,-506719,-506718,-506716,-506715,-506714,-506713,-506712,-506711,-506710,-506709,-506708,-506707,-506706,-506704,-506703,-506702,-506701,-506700,-506699,-506698,-506697,-506696,-506695,-506694,-506692,-506691,-506690,-506689,-506688,-506687,-506686,-506685,-506684,-506683,-506681,-506680,-506679,-506678,-506677,-506676,-506675,-506674,-506673,-506672,-506671,-506669,-506668,-506667,-506666,-506665,-506664,-506663,-506662,-506661,-506660,-506658,-506657,-506656,-506655,-506654,-506653,-506652,-506651,-506650,-506649,-506647,-506646,-506645,-506644,-506643,-506642,-506641,-506640,-506639,-506638,-506636,-506635,-506634,-506633,-506632,-506631,-506630,-506629,-506628,-506627,-506625,-506624,-506623,-506622,-506621,-506620,-506619,-506618,-506617,-506616,-506614,-506613,-506612,-506611,-506610,-506609,-506608,-506607,-506606,-506604,-506603,-506602,-506601,-506600,-506599,-506598,-506597,-506596,-506595,-506593,-506592,-506591,-506590,-506589,-506588,-506587,-506586,-506585,-506583,-506582,-506581,-506580,-506579,-506578,-506577,-506576,-506575,-506573,-506572,-506571,-506570,-506569,-506568,-506567,-506566,-506565,-506564,-506562,-506561,-506560,-506559,-506558,-506557,-506556,-506555,-506554,-506552,-506551,-506550,-506549,-506548,-506547,-506546,-506545,-506544,-506542,-506541,-506540,-506539,-506538,-506537,-506536,-506535,-506533,-506532,-506531,-506530,-506529,-506528,-506527,-506526,-506525,-506523,-506522,-506521,-506520,-506519,-506518,-506517,-506516,-506515,-506513,-506512,-506511,-506510,-506509,-506508,-506507,-506506,-506504,-506503,-506502,-506501,-506500,-506499,-506498,-506497,-506496,-506494,-506493,-506492,-506491,-506490,-506489,-506488,-506487,-506485,-506484,-506483,-506482,-506481,-506480,-506479,-506478,-506477,-506475,-506474,-506473,-506472,-506471,-506470,-506469,-506468,-506466,-506465,-506464,-506463,-506462,-506461,-506460,-506459,-506457,-506456,-506455,-506454,-506453,-506452,-506451,-506450,-506448,-506447,-506446,-506445,-506444,-506443,-506442,-506441,-506439,-506438,-506437,-506436,-506435,-506434,-506433,-506432,-506430,-506429,-506428,-506427,-506426,-506425,-506424,-506423,-506421,-506420,-506419,-506418,-506417,-506416,-506415,-506414,-506412,-506411,-506410,-506409,-506408,-506407,-506406,-506405,-506403,-506402,-506401,-506400,-506399,-506398,-506397,-506396,-506394,-506393,-506392,-506391,-506390,-506389,-506388,-506386,-506385,-506384,-506383,-506382,-506381,-506380,-506379,-506377,-506376,-506375,-506374,-506373,-506372,-506371,-506369,-506368,-506367,-506366,-506365,-506364,-506363,-506362,-506360,-506359,-506358,-506357,-506356,-506355,-506354,-506352,-506351,-506350,-506349,-506348,-506347,-506346,-506345,-506343,-506342,-506341,-506340,-506339,-506338,-506337,-506335,-506334,-506333,-506332,-506331,-506330,-506329,-506327,-506326,-506325,-506324,-506323,-506322,-506321,-506319,-506318,-506317,-506316,-506315,-506314,-506313,-506312,-506310,-506309,-506308,-506307,-506306,-506305,-506304,-506302,-506301,-506300,-506299,-506298,-506297,-506296,-506294,-506293,-506292,-506291,-506290,-506289,-506288,-506286,-506285,-506284,-506283,-506282,-506281,-506280,-506278,-506277,-506276,-506275,-506274,-506273,-506272,-506270,-506269,-506268,-506267,-506266,-506265,-506263,-506262,-506261,-506260,-506259,-506258,-506257,-506255,-506254,-506253,-506252,-506251,-506250,-506249,-506247,-506246,-506245,-506244,-506243,-506242,-506241,-506239,-506238,-506237,-506236,-506235,-506234,-506233,-506231,-506230,-506229,-506228,-506227,-506226,-506224,-506223,-506222,-506221,-506220,-506219,-506218,-506216,-506215,-506214,-506213,-506212,-506211,-506209,-506208,-506207,-506206,-506205,-506204,-506203,-506201,-506200,-506199,-506198,-506197,-506196,-506194,-506193,-506192,-506191,-506190,-506189,-506188,-506186,-506185,-506184,-506183,-506182,-506181,-506179,-506178,-506177,-506176,-506175,-506174,-506173,-506171,-506170,-506169,-506168,-506167,-506166,-506164,-506163,-506162,-506161,-506160,-506159,-506157,-506156,-506155,-506154,-506153,-506152,-506151,-506149,-506148,-506147,-506146,-506145,-506144,-506142,-506141,-506140,-506139,-506138,-506137,-506135,-506134,-506133,-506132,-506131,-506130,-506128,-506127,-506126,-506125,-506124,-506123,-506122,-506120,-506119,-506118,-506117,-506116,-506115,-506113,-506112,-506111,-506110,-506109,-506108,-506106,-506105,-506104,-506103,-506102,-506101,-506099,-506098,-506097,-506096,-506095,-506094,-506092,-506091,-506090,-506089,-506088,-506087,-506085,-506084,-506083,-506082,-506081,-506080,-506078,-506077,-506076,-506075,-506074,-506073,-506071,-506070,-506069,-506068,-506067,-506066,-506064,-506063,-506062,-506061,-506060,-506059,-506057,-506056,-506055,-506054,-506053,-506052,-506050,-506049,-506048,-506047,-506046,-506044,-506043,-506042,-506041,-506040,-506039,-506037,-506036,-506035,-506034,-506033,-506032,-506030,-506029,-506028,-506027,-506026,-506025,-506023,-506022,-506021,-506020,-506019,-506018,-506016,-506015,-506014,-506013,-506012,-506010,-506009,-506008,-506007,-506006,-506005,-506003,-506002,-506001,-506000,-505999,-505998,-505996,-505995,-505994,-505993,-505992,-505990,-505989,-505988,-505987,-505986,-505985,-505983,-505982,-505981,-505980,-505979,-505977,-505976,-505975,-505974,-505973,-505972,-505970,-505969,-505968,-505967,-505966,-505965,-505963,-505962,-505961,-505960,-505959,-505957,-505956,-505955,-505954,-505953,-505952,-505950,-505949,-505948,-505947,-505946,-505944,-505943,-505942,-505941,-505940,-505939,-505937,-505936,-505935,-505934,-505933,-505931,-505930,-505929,-505928,-505927,-505925,-505924,-505923,-505922,-505921,-505920,-505918,-505917,-505916,-505915,-505914,-505912,-505911,-505910,-505909,-505908,-505906,-505905,-505904,-505903,-505902,-505901,-505899,-505898,-505897,-505896,-505895,-505893,-505892,-505891,-505890,-505889,-505887,-505886,-505885,-505884,-505883,-505882,-505880,-505879,-505878,-505877,-505876,-505874,-505873,-505872,-505871,-505870,-505868,-505867,-505866,-505865,-505864,-505862,-505861,-505860,-505859,-505858,-505857,-505855,-505854,-505853,-505852,-505851,-505849,-505848,-505847,-505846,-505845,-505843,-505842,-505841,-505840,-505839,-505837,-505836,-505835,-505834,-505833,-505831,-505830,-505829,-505828,-505827,-505825,-505824,-505823,-505822,-505821,-505819,-505818,-505817,-505816,-505815,-505813,-505812,-505811,-505810,-505809,-505807,-505806,-505805,-505804,-505803,-505801,-505800,-505799,-505798,-505797,-505795,-505794,-505793,-505792,-505791,-505789,-505788,-505787,-505786,-505785,-505783,-505782,-505781,-505780,-505779,-505777,-505776,-505775,-505774,-505773,-505771,-505770,-505769,-505768,-505767,-505765,-505764,-505763,-505762,-505761,-505759,-505758,-505757,-505756,-505755,-505753,-505752,-505751,-505750,-505749,-505747,-505746,-505745,-505744,-505743,-505741,-505740,-505739,-505738,-505737,-505735,-505734,-505733,-505732,-505730,-505729,-505728,-505727,-505726,-505724,-505723,-505722,-505721,-505720,-505718,-505717,-505716,-505715,-505714,-505712,-505711,-505710,-505709,-505708,-505706,-505705,-505704,-505703,-505701,-505700,-505699,-505698,-505697,-505695,-505694,-505693,-505692,-505691,-505689,-505688,-505687,-505686,-505685,-505683,-505682,-505681,-505680,-505678,-505677,-505676,-505675,-505674,-505672,-505671,-505670,-505669,-505668,-505666,-505665,-505664,-505663,-505661,-505660,-505659,-505658,-505657,-505655,-505654,-505653,-505652,-505651,-505649,-505648,-505647,-505646,-505644,-505643,-505642,-505641,-505640,-505638,-505637,-505636,-505635,-505633,-505632,-505631,-505630,-505629,-505627,-505626,-505625,-505624,-505623,-505621,-505620,-505619,-505618,-505616,-505615,-505614,-505613,-505612,-505610,-505609,-505608,-505607,-505605,-505604,-505603,-505602,-505601,-505599,-505598,-505597,-505596,-505594,-505593,-505592,-505591,-505590,-505588,-505587,-505586,-505585,-505583,-505582,-505581,-505580,-505579,-505577,-505576,-505575,-505574,-505572,-505571,-505570,-505569,-505568,-505566,-505565,-505564,-505563,-505561,-505560,-505559,-505558,-505556,-505555,-505554,-505553,-505552,-505550,-505549,-505548,-505547,-505545,-505544,-505543,-505542,-505541,-505539,-505538,-505537,-505536,-505534,-505533,-505532,-505531,-505529,-505528,-505527,-505526,-505525,-505523,-505522,-505521,-505520,-505518,-505517,-505516,-505515,-505513,-505512,-505511,-505510,-505509,-505507,-505506,-505505,-505504,-505502,-505501,-505500,-505499,-505497,-505496,-505495,-505494,-505492,-505491,-505490,-505489,-505488,-505486,-505485,-505484,-505483,-505481,-505480,-505479,-505478,-505476,-505475,-505474,-505473,-505472,-505470,-505469,-505468,-505467,-505465,-505464,-505463,-505462,-505460,-505459,-505458,-505457,-505455,-505454,-505453,-505452,-505450,-505449,-505448,-505447,-505446,-505444,-505443,-505442,-505441,-505439,-505438,-505437,-505436,-505434,-505433,-505432,-505431,-505429,-505428,-505427,-505426,-505424,-505423,-505422,-505421,-505419,-505418,-505417,-505416,-505415,-505413,-505412,-505411,-505410,-505408,-505407,-505406,-505405,-505403,-505402,-505401,-505400,-505398,-505397,-505396,-505395,-505393,-505392,-505391,-505390,-505388,-505387,-505386,-505385,-505383,-505382,-505381,-505380,-505378,-505377,-505376,-505375,-505373,-505372,-505371,-505370,-505368,-505367,-505366,-505365,-505363,-505362,-505361,-505360,-505358,-505357,-505356,-505355,-505353,-505352,-505351,-505350,-505348,-505347,-505346,-505345,-505343,-505342,-505341,-505340,-505338,-505337,-505336,-505335,-505333,-505332,-505331,-505330,-505328,-505327,-505326,-505325,-505323,-505322,-505321,-505320,-505318,-505317,-505316,-505315,-505313,-505312,-505311,-505310,-505308,-505307,-505306,-505305,-505303,-505302,-505301,-505300,-505298,-505297,-505296,-505295,-505293,-505292,-505291,-505290,-505288,-505287,-505286,-505285,-505283,-505282,-505281,-505280,-505278,-505277,-505276,-505275,-505273,-505272,-505271,-505270,-505268,-505267,-505266,-505264,-505263,-505262,-505261,-505259,-505258,-505257,-505256,-505254,-505253,-505252,-505251,-505249,-505248,-505247,-505246,-505244,-505243,-505242,-505241,-505239,-505238,-505237,-505235,-505234,-505233,-505232,-505230,-505229,-505228,-505227,-505225,-505224,-505223,-505222,-505220,-505219,-505218,-505217,-505215,-505214,-505213,-505211,-505210,-505209,-505208,-505206,-505205,-505204,-505203,-505201,-505200,-505199,-505198,-505196,-505195,-505194,-505193,-505191,-505190,-505189,-505187,-505186,-505185,-505184,-505182,-505181,-505180,-505179,-505177,-505176,-505175,-505174,-505172,-505171,-505170,-505168,-505167,-505166,-505165,-505163,-505162,-505161,-505160,-505158,-505157,-505156,-505154,-505153,-505152,-505151,-505149,-505148,-505147,-505146,-505144,-505143,-505142,-505140,-505139,-505138,-505137,-505135,-505134,-505133,-505132,-505130,-505129,-505128,-505126,-505125,-505124,-505123,-505121,-505120,-505119,-505118,-505116,-505115,-505114,-505112,-505111,-505110,-505109,-505107,-505106,-505105,-505104,-505102,-505101,-505100,-505098,-505097,-505096,-505095,-505093,-505092,-505091,-505090,-505088,-505087,-505086,-505084,-505083,-505082,-505081,-505079,-505078,-505077,-505075,-505074,-505073,-505072,-505070,-505069,-505068,-505067,-505065,-505064,-505063,-505061,-505060,-505059,-505058,-505056,-505055,-505054,-505052,-505051,-505050,-505049,-505047,-505046,-505045,-505043,-505042,-505041,-505040,-505038,-505037,-505036,-505034,-505033,-505032,-505031,-505029,-505028,-505027,-505025,-505024,-505023,-505022,-505020,-505019,-505018,-505017,-505015,-505014,-505013,-505011,-505010,-505009,-505008,-505006,-505005,-505004,-505002,-505001,-505000,-504999,-504997,-504996,-504995,-504993,-504992,-504991,-504989,-504988,-504987,-504986,-504984,-504983,-504982,-504980,-504979,-504978,-504977,-504975,-504974,-504973,-504971,-504970,-504969,-504968,-504966,-504965,-504964,-504962,-504961,-504960,-504959,-504957,-504956,-504955,-504953,-504952,-504951,-504950,-504948,-504947,-504946,-504944,-504943,-504942,-504940,-504939,-504938,-504937,-504935,-504934,-504933,-504931,-504930,-504929,-504928,-504926,-504925,-504924,-504922,-504921,-504920,-504918,-504917,-504916,-504915,-504913,-504912,-504911,-504909,-504908,-504907,-504906,-504904,-504903,-504902,-504900,-504899,-504898,-504896,-504895,-504894,-504893,-504891,-504890,-504889,-504887,-504886,-504885,-504883,-504882,-504881,-504880,-504878,-504877,-504876,-504874,-504873,-504872,-504870,-504869,-504868,-504867,-504865,-504864,-504863,-504861,-504860,-504859,-504857,-504856,-504855,-504854,-504852,-504851,-504850,-504848,-504847,-504846,-504844,-504843,-504842,-504841,-504839,-504838,-504837,-504835,-504834,-504833,-504831,-504830,-504829,-504827,-504826,-504825,-504824,-504822,-504821,-504820,-504818,-504817,-504816,-504814,-504813,-504812,-504811,-504809,-504808,-504807,-504805,-504804,-504803,-504801,-504800,-504799,-504797,-504796,-504795,-504794,-504792,-504791,-504790,-504788,-504787,-504786,-504784,-504783,-504782,-504780,-504779,-504778,-504776,-504775,-504774,-504773,-504771,-504770,-504769,-504767,-504766,-504765,-504763,-504762,-504761,-504759,-504758,-504757,-504756,-504754,-504753,-504752,-504750,-504749,-504748,-504746,-504745,-504744,-504742,-504741,-504740,-504738,-504737,-504736,-504735,-504733,-504732,-504731,-504729,-504728,-504727,-504725,-504724,-504723,-504721,-504720,-504719,-504717,-504716,-504715,-504713,-504712,-504711,-504710,-504708,-504707,-504706,-504704,-504703,-504702,-504700,-504699,-504698,-504696,-504695,-504694,-504692,-504691,-504690,-504688,-504687,-504686,-504684,-504683,-504682,-504681,-504679,-504678,-504677,-504675,-504674,-504673,-504671,-504670,-504669,-504667,-504666,-504665,-504663,-504662,-504661,-504659,-504658,-504657,-504655,-504654,-504653,-504651,-504650,-504649,-504647,-504646,-504645,-504644,-504642,-504641,-504640,-504638,-504637,-504636,-504634,-504633,-504632,-504630,-504629,-504628,-504626,-504625,-504624,-504622,-504621,-504620,-504618,-504617,-504616,-504614,-504613,-504612,-504610,-504609,-504608,-504606,-504605,-504604,-504602,-504601,-504600,-504598,-504597,-504596,-504594,-504593,-504592,-504590,-504589,-504588,-504586,-504585,-504584,-504582,-504581,-504580,-504579,-504577,-504576,-504575,-504573,-504572,-504571,-504569,-504568,-504567,-504565,-504564,-504563,-504561,-504560,-504559,-504557,-504556,-504555,-504553,-504552,-504551,-504549,-504548,-504547,-504545,-504544,-504543,-504541,-504540,-504539,-504537,-504536,-504535,-504533,-504532,-504531,-504529,-504528,-504527,-504525,-504524,-504523,-504521,-504520,-504519,-504517,-504516,-504515,-504513,-504512,-504510,-504509,-504508,-504506,-504505,-504504,-504502,-504501,-504500,-504498,-504497,-504496,-504494,-504493,-504492,-504490,-504489,-504488,-504486,-504485,-504484,-504482,-504481,-504480,-504478,-504477,-504476,-504474,-504473,-504472,-504470,-504469,-504468,-504466,-504465,-504464,-504462,-504461,-504460,-504458,-504457,-504456,-504454,-504453,-504452,-504450,-504449,-504448,-504446,-504445,-504443,-504442,-504441,-504439,-504438,-504437,-504435,-504434,-504433,-504431,-504430,-504429,-504427,-504426,-504425,-504423,-504422,-504421,-504419,-504418,-504417,-504415,-504414,-504413,-504411,-504410,-504408,-504407,-504406,-504404,-504403,-504402,-504400,-504399,-504398,-504396,-504395,-504394,-504392,-504391,-504390,-504388,-504387,-504386,-504384,-504383,-504382,-504380,-504379,-504377,-504376,-504375,-504373,-504372,-504371,-504369,-504368,-504367,-504365,-504364,-504363,-504361,-504360,-504359,-504357,-504356,-504354,-504353,-504352,-504350,-504349,-504348,-504346,-504345,-504344,-504342,-504341,-504340,-504338,-504337,-504336,-504334,-504333,-504331,-504330,-504329,-504327,-504326,-504325,-504323,-504322,-504321,-504319,-504318,-504317,-504315,-504314,-504312,-504311,-504310,-504308,-504307,-504306,-504304,-504303,-504302,-504300,-504299,-504298,-504296,-504295,-504293,-504292,-504291,-504289,-504288,-504287,-504285,-504284,-504283,-504281,-504280,-504279,-504277,-504276,-504274,-504273,-504272,-504270,-504269,-504268,-504266,-504265,-504264,-504262,-504261,-504259,-504258,-504257,-504255,-504254,-504253,-504251,-504250,-504249,-504247,-504246,-504244,-504243,-504242,-504240,-504239,-504238,-504236,-504235,-504234,-504232,-504231,-504229,-504228,-504227,-504225,-504224,-504223,-504221,-504220,-504219,-504217,-504216,-504214,-504213,-504212,-504210,-504209,-504208,-504206,-504205,-504204,-504202,-504201,-504199,-504198,-504197,-504195,-504194,-504193,-504191,-504190,-504188,-504187,-504186,-504184,-504183,-504182,-504180,-504179,-504178,-504176,-504175,-504173,-504172,-504171,-504169,-504168,-504167,-504165,-504164,-504162,-504161,-504160,-504158,-504157,-504156,-504154,-504153,-504151,-504150,-504149,-504147,-504146,-504145,-504143,-504142,-504140,-504139,-504138,-504136,-504135,-504134,-504132,-504131,-504129,-504128,-504127,-504125,-504124,-504123,-504121,-504120,-504118,-504117,-504116,-504114,-504113,-504112,-504110,-504109,-504107,-504106,-504105,-504103,-504102,-504101,-504099,-504098,-504096,-504095,-504094,-504092,-504091,-504090,-504088,-504087,-504085,-504084,-504083,-504081,-504080,-504079,-504077,-504076,-504074,-504073,-504072,-504070,-504069,-504067,-504066,-504065,-504063,-504062,-504061,-504059,-504058,-504056,-504055,-504054,-504052,-504051,-504049,-504048,-504047,-504045,-504044,-504043,-504041,-504040,-504038,-504037,-504036,-504034,-504033,-504032,-504030,-504029,-504027,-504026,-504025,-504023,-504022,-504020,-504019,-504018,-504016,-504015,-504014,-504012,-504011,-504009,-504008,-504007,-504005,-504004,-504002,-504001,-504000,-503998,-503997,-503995,-503994,-503993,-503991,-503990,-503989,-503987,-503986,-503984,-503983,-503982,-503980,-503979,-503977,-503976,-503975,-503973,-503972,-503970,-503969,-503968,-503966,-503965,-503964,-503962,-503961,-503959,-503958,-503957,-503955,-503954,-503952,-503951,-503950,-503948,-503947,-503945,-503944,-503943,-503941,-503940,-503938,-503937,-503936,-503934,-503933,-503931,-503930,-503929,-503927,-503926,-503925,-503923,-503922,-503920,-503919,-503918,-503916,-503915,-503913,-503912,-503911,-503909,-503908,-503906,-503905,-503904,-503902,-503901,-503899,-503898,-503897,-503895,-503894,-503892,-503891,-503890,-503888,-503887,-503885,-503884,-503883,-503881,-503880,-503878,-503877,-503876,-503874,-503873,-503871,-503870,-503869,-503867,-503866,-503864,-503863,-503862,-503860,-503859,-503857,-503856,-503855,-503853,-503852,-503850,-503849,-503848,-503846,-503845,-503843,-503842,-503841,-503839,-503838,-503836,-503835,-503834,-503832,-503831,-503829,-503828,-503827,-503825,-503824,-503822,-503821,-503820,-503818,-503817,-503815,-503814,-503812,-503811,-503810,-503808,-503807,-503805,-503804,-503803,-503801,-503800,-503798,-503797,-503796,-503794,-503793,-503791,-503790,-503789,-503787,-503786,-503784,-503783,-503782,-503780,-503779,-503777,-503776,-503774,-503773,-503772,-503770,-503769,-503767,-503766,-503765,-503763,-503762,-503760,-503759,-503758,-503756,-503755,-503753,-503752,-503751,-503749,-503748,-503746,-503745,-503743,-503742,-503741,-503739,-503738,-503736,-503735,-503734,-503732,-503731,-503729,-503728,-503726,-503725,-503724,-503722,-503721,-503719,-503718,-503717,-503715,-503714,-503712,-503711,-503710,-503708,-503707,-503705,-503704,-503702,-503701,-503700,-503698,-503697,-503695,-503694,-503693,-503691,-503690,-503688,-503687,-503685,-503684,-503683,-503681,-503680,-503678,-503677,-503675,-503674,-503673,-503671,-503670,-503668,-503667,-503666,-503664,-503663,-503661,-503660,-503658,-503657,-503656,-503654,-503653,-503651,-503650,-503649,-503647,-503646,-503644,-503643,-503641,-503640,-503639,-503637,-503636,-503634,-503633,-503631,-503630,-503629,-503627,-503626,-503624,-503623,-503621,-503620,-503619,-503617,-503616,-503614,-503613,-503612,-503610,-503609,-503607,-503606,-503604,-503603,-503602,-503600,-503599,-503597,-503596,-503594,-503593,-503592,-503590,-503589,-503587,-503586,-503584,-503583,-503582,-503580,-503579,-503577,-503576,-503574,-503573,-503572,-503570,-503569,-503567,-503566,-503564,-503563,-503562,-503560,-503559,-503557,-503556,-503554,-503553,-503552,-503550,-503549,-503547,-503546,-503544,-503543,-503542,-503540,-503539,-503537,-503536,-503534,-503533,-503532,-503530,-503529,-503527,-503526,-503524,-503523,-503521,-503520,-503519,-503517,-503516,-503514,-503513,-503511,-503510,-503509,-503507,-503506,-503504,-503503,-503501,-503500,-503499,-503497,-503496,-503494,-503493,-503491,-503490,-503488,-503487,-503486,-503484,-503483,-503481,-503480,-503478,-503477,-503476,-503474,-503473,-503471,-503470,-503468,-503467,-503465,-503464,-503463,-503461,-503460,-503458,-503457,-503455,-503454,-503453,-503451,-503450,-503448,-503447,-503445,-503444,-503442,-503441,-503440,-503438,-503437,-503435,-503434,-503432,-503431,-503429,-503428,-503427,-503425,-503424,-503422,-503421,-503419,-503418,-503416,-503415,-503414,-503412,-503411,-503409,-503408,-503406,-503405,-503403,-503402,-503401,-503399,-503398,-503396,-503395,-503393,-503392,-503390,-503389,-503388,-503386,-503385,-503383,-503382,-503380,-503379,-503377,-503376,-503375,-503373,-503372,-503370,-503369,-503367,-503366,-503364,-503363,-503362,-503360,-503359,-503357,-503356,-503354,-503353,-503351,-503350,-503349,-503347,-503346,-503344,-503343,-503341,-503340,-503338,-503337,-503335,-503334,-503333,-503331,-503330,-503328,-503327,-503325,-503324,-503322,-503321,-503319,-503318,-503317,-503315,-503314,-503312,-503311,-503309,-503308,-503306,-503305,-503304,-503302,-503301,-503299,-503298,-503296,-503295,-503293,-503292,-503290,-503289,-503288,-503286,-503285,-503283,-503282,-503280,-503279,-503277,-503276,-503274,-503273,-503272,-503270,-503269,-503267,-503266,-503264,-503263,-503261,-503260,-503258,-503257,-503255,-503254,-503253,-503251,-503250,-503248,-503247,-503245,-503244,-503242,-503241,-503239,-503238,-503237,-503235,-503234,-503232,-503231,-503229,-503228,-503226,-503225,-503223,-503222,-503220,-503219,-503218,-503216,-503215,-503213,-503212,-503210,-503209,-503207,-503206,-503204,-503203,-503201,-503200,-503199,-503197,-503196,-503194,-503193,-503191,-503190,-503188,-503187,-503185,-503184,-503182,-503181,-503179,-503178,-503177,-503175,-503174,-503172,-503171,-503169,-503168,-503166,-503165,-503163,-503162,-503160,-503159,-503157,-503156,-503155,-503153,-503152,-503150,-503149,-503147,-503146,-503144,-503143,-503141,-503140,-503138,-503137,-503135,-503134,-503133,-503131,-503130,-503128,-503127,-503125,-503124,-503122,-503121,-503119,-503118,-503116,-503115,-503113,-503112,-503110,-503109,-503108,-503106,-503105,-503103,-503102,-503100,-503099,-503097,-503096,-503094,-503093,-503091,-503090,-503088,-503087,-503085,-503084,-503082,-503081,-503080,-503078,-503077,-503075,-503074,-503072,-503071,-503069,-503068,-503066,-503065,-503063,-503062,-503060,-503059,-503057,-503056,-503054,-503053,-503051,-503050,-503049,-503047,-503046,-503044,-503043,-503041,-503040,-503038,-503037,-503035,-503034,-503032,-503031,-503029,-503028,-503026,-503025,-503023,-503022,-503020,-503019,-503017,-503016,-503015,-503013,-503012,-503010,-503009,-503007,-503006,-503004,-503003,-503001,-503000,-502998,-502997,-502995,-502994,-502992,-502991,-502989,-502988,-502986,-502985,-502983,-502982,-502980,-502979,-502977,-502976,-502975,-502973,-502972,-502970,-502969,-502967,-502966,-502964,-502963,-502961,-502960,-502958,-502957,-502955,-502954,-502952,-502951,-502949,-502948,-502946,-502945,-502943,-502942,-502940,-502939,-502937,-502936,-502934,-502933,-502931,-502930,-502928,-502927,-502925,-502924,-502922,-502921,-502920,-502918,-502917,-502915,-502914,-502912,-502911,-502909,-502908,-502906,-502905,-502903,-502902,-502900,-502899,-502897,-502896,-502894,-502893,-502891,-502890,-502888,-502887,-502885,-502884,-502882,-502881,-502879,-502878,-502876,-502875,-502873,-502872,-502870,-502869,-502867,-502866,-502864,-502863,-502861,-502860,-502858,-502857,-502855,-502854,-502852,-502851,-502849,-502848,-502846,-502845,-502843,-502842,-502840,-502839,-502837,-502836,-502834,-502833,-502831,-502830,-502828,-502827,-502825,-502824,-502822,-502821,-502819,-502818,-502816,-502815,-502813,-502812,-502810,-502809,-502807,-502806,-502804,-502803,-502801,-502800,-502798,-502797,-502795,-502794,-502792,-502791,-502789,-502788,-502786,-502785,-502783,-502782,-502780,-502779,-502777,-502776,-502774,-502773,-502771,-502770,-502768,-502767,-502765,-502764,-502762,-502761,-502759,-502758,-502756,-502755,-502753,-502752,-502750,-502749,-502747,-502746,-502744,-502743,-502741,-502740,-502738,-502737,-502735,-502734,-502732,-502731,-502729,-502728,-502726,-502725,-502723,-502722,-502720,-502719,-502717,-502716,-502714,-502713,-502711,-502710,-502708,-502707,-502705,-502704,-502702,-502701,-502699,-502698,-502696,-502695,-502693,-502692,-502690,-502689,-502687,-502686,-502684,-502683,-502681,-502680,-502678,-502677,-502675,-502674,-502672,-502671,-502669,-502667,-502666,-502664,-502663,-502661,-502660,-502658,-502657,-502655,-502654,-502652,-502651,-502649,-502648,-502646,-502645,-502643,-502642,-502640,-502639,-502637,-502636,-502634,-502633,-502631,-502630,-502628,-502627,-502625,-502624,-502622,-502621,-502619,-502618,-502616,-502615,-502613,-502611,-502610,-502608,-502607,-502605,-502604,-502602,-502601,-502599,-502598,-502596,-502595,-502593,-502592,-502590,-502589,-502587,-502586,-502584,-502583,-502581,-502580,-502578,-502577,-502575,-502574,-502572,-502570,-502569,-502567,-502566,-502564,-502563,-502561,-502560,-502558,-502557,-502555,-502554,-502552,-502551,-502549,-502548,-502546,-502545,-502543,-502542,-502540,-502539,-502537,-502535,-502534,-502532,-502531,-502529,-502528,-502526,-502525,-502523,-502522,-502520,-502519,-502517,-502516,-502514,-502513,-502511,-502510,-502508,-502507,-502505,-502503,-502502,-502500,-502499,-502497,-502496,-502494,-502493,-502491,-502490,-502488,-502487,-502485,-502484,-502482,-502481,-502479,-502478,-502476,-502474,-502473,-502471,-502470,-502468,-502467,-502465,-502464,-502462,-502461,-502459,-502458,-502456,-502455,-502453,-502452,-502450,-502448,-502447,-502445,-502444,-502442,-502441,-502439,-502438,-502436,-502435,-502433,-502432,-502430,-502429,-502427,-502425,-502424,-502422,-502421,-502419,-502418,-502416,-502415,-502413,-502412,-502410,-502409,-502407,-502406,-502404,-502402,-502401,-502399,-502398,-502396,-502395,-502393,-502392,-502390,-502389,-502387,-502386,-502384,-502382,-502381,-502379,-502378,-502376,-502375,-502373,-502372,-502370,-502369,-502367,-502366,-502364,-502363,-502361,-502359,-502358,-502356,-502355,-502353,-502352,-502350,-502349,-502347,-502346,-502344,-502343,-502341,-502339,-502338,-502336,-502335,-502333,-502332,-502330,-502329,-502327,-502326,-502324,-502322,-502321,-502319,-502318,-502316,-502315,-502313,-502312,-502310,-502309,-502307,-502306,-502304,-502302,-502301,-502299,-502298,-502296,-502295,-502293,-502292,-502290,-502289,-502287,-502285,-502284,-502282,-502281,-502279,-502278,-502276,-502275,-502273,-502272,-502270,-502268,-502267,-502265,-502264,-502262,-502261,-502259,-502258,-502256,-502254,-502253,-502251,-502250,-502248,-502247,-502245,-502244,-502242,-502241,-502239,-502237,-502236,-502234,-502233,-502231,-502230,-502228,-502227,-502225,-502224,-502222,-502220,-502219,-502217,-502216,-502214,-502213,-502211,-502210,-502208,-502206,-502205,-502203,-502202,-502200,-502199,-502197,-502196,-502194,-502192,-502191,-502189,-502188,-502186,-502185,-502183,-502182,-502180,-502178,-502177,-502175,-502174,-502172,-502171,-502169,-502168,-502166,-502165,-502163,-502161,-502160,-502158,-502157,-502155,-502154,-502152,-502150,-502149,-502147,-502146,-502144,-502143,-502141,-502140,-502138,-502136,-502135,-502133,-502132,-502130,-502129,-502127,-502126,-502124,-502122,-502121,-502119,-502118,-502116,-502115,-502113,-502112,-502110,-502108,-502107,-502105,-502104,-502102,-502101,-502099,-502097,-502096,-502094,-502093,-502091,-502090,-502088,-502087,-502085,-502083,-502082,-502080,-502079,-502077,-502076,-502074,-502072,-502071,-502069,-502068,-502066,-502065,-502063,-502062,-502060,-502058,-502057,-502055,-502054,-502052,-502051,-502049,-502047,-502046,-502044,-502043,-502041,-502040,-502038,-502036,-502035,-502033,-502032,-502030,-502029,-502027,-502026,-502024,-502022,-502021,-502019,-502018,-502016,-502015,-502013,-502011,-502010,-502008,-502007,-502005,-502004,-502002,-502000,-501999,-501997,-501996,-501994,-501993,-501991,-501989,-501988,-501986,-501985,-501983,-501982,-501980,-501978,-501977,-501975,-501974,-501972,-501971,-501969,-501967,-501966,-501964,-501963,-501961,-501960,-501958,-501956,-501955,-501953,-501952,-501950,-501949,-501947,-501945,-501944,-501942,-501941,-501939,-501938,-501936,-501934,-501933,-501931,-501930,-501928,-501927,-501925,-501923,-501922,-501920,-501919,-501917,-501915,-501914,-501912,-501911,-501909,-501908,-501906,-501904,-501903,-501901,-501900,-501898,-501897,-501895,-501893,-501892,-501890,-501889,-501887,-501885,-501884,-501882,-501881,-501879,-501878,-501876,-501874,-501873,-501871,-501870,-501868,-501867,-501865,-501863,-501862,-501860,-501859,-501857,-501855,-501854,-501852,-501851,-501849,-501848,-501846,-501844,-501843,-501841,-501840,-501838,-501836,-501835,-501833,-501832,-501830,-501829,-501827,-501825,-501824,-501822,-501821,-501819,-501817,-501816,-501814,-501813,-501811,-501810,-501808,-501806,-501805,-501803,-501802,-501800,-501798,-501797,-501795,-501794,-501792,-501790,-501789,-501787,-501786,-501784,-501783,-501781,-501779,-501778,-501776,-501775,-501773,-501771,-501770,-501768,-501767,-501765,-501763,-501762,-501760,-501759,-501757,-501756,-501754,-501752,-501751,-501749,-501748,-501746,-501744,-501743,-501741,-501740,-501738,-501736,-501735,-501733,-501732,-501730,-501728,-501727,-501725,-501724,-501722,-501720,-501719,-501717,-501716,-501714,-501713,-501711,-501709,-501708,-501706,-501705,-501703,-501701,-501700,-501698,-501697,-501695,-501693,-501692,-501690,-501689,-501687,-501685,-501684,-501682,-501681,-501679,-501677,-501676,-501674,-501673,-501671,-501669,-501668,-501666,-501665,-501663,-501661,-501660,-501658,-501657,-501655,-501653,-501652,-501650,-501649,-501647,-501645,-501644,-501642,-501641,-501639,-501637,-501636,-501634,-501633,-501631,-501629,-501628,-501626,-501625,-501623,-501621,-501620,-501618,-501617,-501615,-501613,-501612,-501610,-501609,-501607,-501605,-501604,-501602,-501601,-501599,-501597,-501596,-501594,-501593,-501591,-501589,-501588,-501586,-501585,-501583,-501581,-501580,-501578,-501577,-501575,-501573,-501572,-501570,-501569,-501567,-501565,-501564,-501562,-501560,-501559,-501557,-501556,-501554,-501552,-501551,-501549,-501548,-501546,-501544,-501543,-501541,-501540,-501538,-501536,-501535,-501533,-501532,-501530,-501528,-501527,-501525,-501523,-501522,-501520,-501519,-501517,-501515,-501514,-501512,-501511,-501509,-501507,-501506,-501504,-501503,-501501,-501499,-501498,-501496,-501494,-501493,-501491,-501490,-501488,-501486,-501485,-501483,-501482,-501480,-501478,-501477,-501475,-501473,-501472,-501470,-501469,-501467,-501465,-501464,-501462,-501461,-501459,-501457,-501456,-501454,-501453,-501451,-501449,-501448,-501446,-501444,-501443,-501441,-501440,-501438,-501436,-501435,-501433,-501431,-501430,-501428,-501427,-501425,-501423,-501422,-501420,-501419,-501417,-501415,-501414,-501412,-501410,-501409,-501407,-501406,-501404,-501402,-501401,-501399,-501397,-501396,-501394,-501393,-501391,-501389,-501388,-501386,-501385,-501383,-501381,-501380,-501378,-501376,-501375,-501373,-501372,-501370,-501368,-501367,-501365,-501363,-501362,-501360,-501359,-501357,-501355,-501354,-501352,-501350,-501349,-501347,-501346,-501344,-501342,-501341,-501339,-501337,-501336,-501334,-501333,-501331,-501329,-501328,-501326,-501324,-501323,-501321,-501320,-501318,-501316,-501315,-501313,-501311,-501310,-501308,-501307,-501305,-501303,-501302,-501300,-501298,-501297,-501295,-501294,-501292,-501290,-501289,-501287,-501285,-501284,-501282,-501280,-501279,-501277,-501276,-501274,-501272,-501271,-501269,-501267,-501266,-501264,-501263,-501261,-501259,-501258,-501256,-501254,-501253,-501251,-501249,-501248,-501246,-501245,-501243,-501241,-501240,-501238,-501236,-501235,-501233,-501232,-501230,-501228,-501227,-501225,-501223,-501222,-501220,-501218,-501217,-501215,-501214,-501212,-501210,-501209,-501207,-501205,-501204,-501202,-501200,-501199,-501197,-501196,-501194,-501192,-501191,-501189,-501187,-501186,-501184,-501182,-501181,-501179,-501178,-501176,-501174,-501173,-501171,-501169,-501168,-501166,-501164,-501163,-501161,-501159,-501158,-501156,-501155,-501153,-501151,-501150,-501148,-501146,-501145,-501143,-501141,-501140,-501138,-501136,-501135,-501133,-501132,-501130,-501128,-501127,-501125,-501123,-501122,-501120,-501118,-501117,-501115,-501113,-501112,-501110,-501109,-501107,-501105,-501104,-501102,-501100,-501099,-501097,-501095,-501094,-501092,-501090,-501089,-501087,-501086,-501084,-501082,-501081,-501079,-501077,-501076,-501074,-501072,-501071,-501069,-501067,-501066,-501064,-501062,-501061,-501059,-501058,-501056,-501054,-501053,-501051,-501049,-501048,-501046,-501044,-501043,-501041,-501039,-501038,-501036,-501034,-501033,-501031,-501029,-501028,-501026,-501025,-501023,-501021,-501020,-501018,-501016,-501015,-501013,-501011,-501010,-501008,-501006,-501005,-501003,-501001,-501000,-500998,-500996,-500995,-500993,-500991,-500990,-500988,-500987,-500985,-500983,-500982,-500980,-500978,-500977,-500975,-500973,-500972,-500970,-500968,-500967,-500965,-500963,-500962,-500960,-500958,-500957,-500955,-500953,-500952,-500950,-500948,-500947,-500945,-500943,-500942,-500940,-500938,-500937,-500935,-500934,-500932,-500930,-500929,-500927,-500925,-500924,-500922,-500920,-500919,-500917,-500915,-500914,-500912,-500910,-500909,-500907,-500905,-500904,-500902,-500900,-500899,-500897,-500895,-500894,-500892,-500890,-500889,-500887,-500885,-500884,-500882,-500880,-500879,-500877,-500875,-500874,-500872,-500870,-500869,-500867,-500865,-500864,-500862,-500860,-500859,-500857,-500855,-500854,-500852,-500850,-500849,-500847,-500845,-500844,-500842,-500840,-500839,-500837,-500835,-500834,-500832,-500830,-500829,-500827,-500825,-500824,-500822,-500820,-500819,-500817,-500815,-500814,-500812,-500810,-500809,-500807,-500805,-500804,-500802,-500800,-500799,-500797,-500795,-500794,-500792,-500790,-500789,-500787,-500785,-500784,-500782,-500780,-500779,-500777,-500775,-500774,-500772,-500770,-500769,-500767,-500765,-500764,-500762,-500760,-500759,-500757,-500755,-500754,-500752,-500750,-500749,-500747,-500745,-500744,-500742,-500740,-500739,-500737,-500735,-500734,-500732,-500730,-500729,-500727,-500725,-500723,-500722,-500720,-500718,-500717,-500715,-500713,-500712,-500710,-500708,-500707,-500705,-500703,-500702,-500700,-500698,-500697,-500695,-500693,-500692,-500690,-500688,-500687,-500685,-500683,-500682,-500680,-500678,-500677,-500675,-500673,-500671,-500670,-500668,-500666,-500665,-500663,-500661,-500660,-500658,-500656,-500655,-500653,-500651,-500650,-500648,-500646,-500645,-500643,-500641,-500640,-500638,-500636,-500635,-500633,-500631,-500629,-500628,-500626,-500624,-500623,-500621,-500619,-500618,-500616,-500614,-500613,-500611,-500609,-500608,-500606,-500604,-500603,-500601,-500599,-500597,-500596,-500594,-500592,-500591,-500589,-500587,-500586,-500584,-500582,-500581,-500579,-500577,-500576,-500574,-500572,-500570,-500569,-500567,-500565,-500564,-500562,-500560,-500559,-500557,-500555,-500554,-500552,-500550,-500549,-500547,-500545,-500543,-500542,-500540,-500538,-500537,-500535,-500533,-500532,-500530,-500528,-500527,-500525,-500523,-500521,-500520,-500518,-500516,-500515,-500513,-500511,-500510,-500508,-500506,-500505,-500503,-500501,-500499,-500498,-500496,-500494,-500493,-500491,-500489,-500488,-500486,-500484,-500483,-500481,-500479,-500477,-500476,-500474,-500472,-500471,-500469,-500467,-500466,-500464,-500462,-500461,-500459,-500457,-500455,-500454,-500452,-500450,-500449,-500447,-500445,-500444,-500442,-500440,-500438,-500437,-500435,-500433,-500432,-500430,-500428,-500427,-500425,-500423,-500421,-500420,-500418,-500416,-500415,-500413,-500411,-500410,-500408,-500406,-500404,-500403,-500401,-500399,-500398,-500396,-500394,-500393,-500391,-500389,-500387,-500386,-500384,-500382,-500381,-500379,-500377,-500376,-500374,-500372,-500370,-500369,-500367,-500365,-500364,-500362,-500360,-500359,-500357,-500355,-500353,-500352,-500350,-500348,-500347,-500345,-500343,-500341,-500340,-500338,-500336,-500335,-500333,-500331,-500330,-500328,-500326,-500324,-500323,-500321,-500319,-500318,-500316,-500314,-500312,-500311,-500309,-500307,-500306,-500304,-500302,-500300,-500299,-500297,-500295,-500294,-500292,-500290,-500289,-500287,-500285,-500283,-500282,-500280,-500278,-500277,-500275,-500273,-500271,-500270,-500268,-500266,-500265,-500263,-500261,-500259,-500258,-500256,-500254,-500253,-500251,-500249,-500247,-500246,-500244,-500242,-500241,-500239,-500237,-500235,-500234,-500232,-500230,-500229,-500227,-500225,-500223,-500222,-500220,-500218,-500217,-500215,-500213,-500211,-500210,-500208,-500206,-500205,-500203,-500201,-500199,-500198,-500196,-500194,-500193,-500191,-500189,-500187,-500186,-500184,-500182,-500181,-500179,-500177,-500175,-500174,-500172,-500170,-500169,-500167,-500165,-500163,-500162,-500160,-500158,-500156,-500155,-500153,-500151,-500150,-500148,-500146,-500144,-500143,-500141,-500139,-500138,-500136,-500134,-500132,-500131,-500129,-500127,-500125,-500124,-500122,-500120,-500119,-500117,-500115,-500113,-500112,-500110,-500108,-500107,-500105,-500103,-500101,-500100,-500098,-500096,-500094,-500093,-500091,-500089,-500088,-500086,-500084,-500082,-500081,-500079,-500077,-500075,-500074,-500072,-500070,-500069,-500067,-500065,-500063,-500062,-500060,-500058,-500056,-500055,-500053,-500051,-500050,-500048,-500046,-500044,-500043,-500041,-500039,-500037,-500036,-500034,-500032,-500031,-500029,-500027,-500025,-500024,-500022,-500020,-500018,-500017,-500015,-500013,-500012,-500010,-500008,-500006,-500005,-500003,-500001,-499999,-499998,-499996,-499994,-499992,-499991,-499989,-499987,-499986,-499984,-499982,-499980,-499979,-499977,-499975,-499973,-499972,-499970,-499968,-499966,-499965,-499963,-499961,-499960,-499958,-499956,-499954,-499953,-499951,-499949,-499947,-499946,-499944,-499942,-499940,-499939,-499937,-499935,-499933,-499932,-499930,-499928,-499927,-499925,-499923,-499921,-499920,-499918,-499916,-499914,-499913,-499911,-499909,-499907,-499906,-499904,-499902,-499900,-499899,-499897,-499895,-499893,-499892,-499890,-499888,-499887,-499885,-499883,-499881,-499880,-499878,-499876,-499874,-499873,-499871,-499869,-499867,-499866,-499864,-499862,-499860,-499859,-499857,-499855,-499853,-499852,-499850,-499848,-499846,-499845,-499843,-499841,-499839,-499838,-499836,-499834,-499832,-499831,-499829,-499827,-499825,-499824,-499822,-499820,-499819,-499817,-499815,-499813,-499812,-499810,-499808,-499806,-499805,-499803,-499801,-499799,-499798,-499796,-499794,-499792,-499791,-499789,-499787,-499785,-499784,-499782,-499780,-499778,-499777,-499775,-499773,-499771,-499770,-499768,-499766,-499764,-499763,-499761,-499759,-499757,-499756,-499754,-499752,-499750,-499749,-499747,-499745,-499743,-499742,-499740,-499738,-499736,-499735,-499733,-499731,-499729,-499728,-499726,-499724,-499722,-499721,-499719,-499717,-499715,-499713,-499712,-499710,-499708,-499706,-499705,-499703,-499701,-499699,-499698,-499696,-499694,-499692,-499691,-499689,-499687,-499685,-499684,-499682,-499680,-499678,-499677,-499675,-499673,-499671,-499670,-499668,-499666,-499664,-499663,-499661,-499659,-499657,-499656,-499654,-499652,-499650,-499648,-499647,-499645,-499643,-499641,-499640,-499638,-499636,-499634,-499633,-499631,-499629,-499627,-499626,-499624,-499622,-499620,-499619,-499617,-499615,-499613,-499612,-499610,-499608,-499606,-499604,-499603,-499601,-499599,-499597,-499596,-499594,-499592,-499590,-499589,-499587,-499585,-499583,-499582,-499580,-499578,-499576,-499574,-499573,-499571,-499569,-499567,-499566,-499564,-499562,-499560,-499559,-499557,-499555,-499553,-499552,-499550,-499548,-499546,-499544,-499543,-499541,-499539,-499537,-499536,-499534,-499532,-499530,-499529,-499527,-499525,-499523,-499521,-499520,-499518,-499516,-499514,-499513,-499511,-499509,-499507,-499506,-499504,-499502,-499500,-499498,-499497,-499495,-499493,-499491,-499490,-499488,-499486,-499484,-499483,-499481,-499479,-499477,-499475,-499474,-499472,-499470,-499468,-499467,-499465,-499463,-499461,-499460,-499458,-499456,-499454,-499452,-499451,-499449,-499447,-499445,-499444,-499442,-499440,-499438,-499436,-499435,-499433,-499431,-499429,-499428,-499426,-499424,-499422,-499420,-499419,-499417,-499415,-499413,-499412,-499410,-499408,-499406,-499404,-499403,-499401,-499399,-499397,-499396,-499394,-499392,-499390,-499388,-499387,-499385,-499383,-499381,-499380,-499378,-499376,-499374,-499372,-499371,-499369,-499367,-499365,-499364,-499362,-499360,-499358,-499356,-499355,-499353,-499351,-499349,-499348,-499346,-499344,-499342,-499340,-499339,-499337,-499335,-499333,-499331,-499330,-499328,-499326,-499324,-499323,-499321,-499319,-499317,-499315,-499314,-499312,-499310,-499308,-499306,-499305,-499303,-499301,-499299,-499298,-499296,-499294,-499292,-499290,-499289,-499287,-499285,-499283,-499281,-499280,-499278,-499276,-499274,-499273,-499271,-499269,-499267,-499265,-499264,-499262,-499260,-499258,-499256,-499255,-499253,-499251,-499249,-499248,-499246,-499244,-499242,-499240,-499239,-499237,-499235,-499233,-499231,-499230,-499228,-499226,-499224,-499222,-499221,-499219,-499217,-499215,-499213,-499212,-499210,-499208,-499206,-499205,-499203,-499201,-499199,-499197,-499196,-499194,-499192,-499190,-499188,-499187,-499185,-499183,-499181,-499179,-499178,-499176,-499174,-499172,-499170,-499169,-499167,-499165,-499163,-499161,-499160,-499158,-499156,-499154,-499152,-499151,-499149,-499147,-499145,-499144,-499142,-499140,-499138,-499136,-499135,-499133,-499131,-499129,-499127,-499126,-499124,-499122,-499120,-499118,-499117,-499115,-499113,-499111,-499109,-499108,-499106,-499104,-499102,-499100,-499099,-499097,-499095,-499093,-499091,-499090,-499088,-499086,-499084,-499082,-499081,-499079,-499077,-499075,-499073,-499072,-499070,-499068,-499066,-499064,-499062,-499061,-499059,-499057,-499055,-499053,-499052,-499050,-499048,-499046,-499044,-499043,-499041,-499039,-499037,-499035,-499034,-499032,-499030,-499028,-499026,-499025,-499023,-499021,-499019,-499017,-499016,-499014,-499012,-499010,-499008,-499007,-499005,-499003,-499001,-498999,-498997,-498996,-498994,-498992,-498990,-498988,-498987,-498985,-498983,-498981,-498979,-498978,-498976,-498974,-498972,-498970,-498969,-498967,-498965,-498963,-498961,-498960,-498958,-498956,-498954,-498952,-498950,-498949,-498947,-498945,-498943,-498941,-498940,-498938,-498936,-498934,-498932,-498931,-498929,-498927,-498925,-498923,-498921,-498920,-498918,-498916,-498914,-498912,-498911,-498909,-498907,-498905,-498903,-498901,-498900,-498898,-498896,-498894,-498892,-498891,-498889,-498887,-498885,-498883,-498882,-498880,-498878,-498876,-498874,-498872,-498871,-498869,-498867,-498865,-498863,-498862,-498860,-498858,-498856,-498854,-498852,-498851,-498849,-498847,-498845,-498843,-498842,-498840,-498838,-498836,-498834,-498832,-498831,-498829,-498827,-498825,-498823,-498821,-498820,-498818,-498816,-498814,-498812,-498811,-498809,-498807,-498805,-498803,-498801,-498800,-498798,-498796,-498794,-498792,-498791,-498789,-498787,-498785,-498783,-498781,-498780,-498778,-498776,-498774,-498772,-498770,-498769,-498767,-498765,-498763,-498761,-498760,-498758,-498756,-498754,-498752,-498750,-498749,-498747,-498745,-498743,-498741,-498739,-498738,-498736,-498734,-498732,-498730,-498728,-498727,-498725,-498723,-498721,-498719,-498717,-498716,-498714,-498712,-498710,-498708,-498707,-498705,-498703,-498701,-498699,-498697,-498696,-498694,-498692,-498690,-498688,-498686,-498685,-498683,-498681,-498679,-498677,-498675,-498674,-498672,-498670,-498668,-498666,-498664,-498663,-498661,-498659,-498657,-498655,-498653,-498652,-498650,-498648,-498646,-498644,-498642,-498641,-498639,-498637,-498635,-498633,-498631,-498630,-498628,-498626,-498624,-498622,-498620,-498619,-498617,-498615,-498613,-498611,-498609,-498608,-498606,-498604,-498602,-498600,-498598,-498597,-498595,-498593,-498591,-498589,-498587,-498585,-498584,-498582,-498580,-498578,-498576,-498574,-498573,-498571,-498569,-498567,-498565,-498563,-498562,-498560,-498558,-498556,-498554,-498552,-498551,-498549,-498547,-498545,-498543,-498541,-498539,-498538,-498536,-498534,-498532,-498530,-498528,-498527,-498525,-498523,-498521,-498519,-498517,-498516,-498514,-498512,-498510,-498508,-498506,-498504,-498503,-498501,-498499,-498497,-498495,-498493,-498492,-498490,-498488,-498486,-498484,-498482,-498480,-498479,-498477,-498475,-498473,-498471,-498469,-498468,-498466,-498464,-498462,-498460,-498458,-498456,-498455,-498453,-498451,-498449,-498447,-498445,-498444,-498442,-498440,-498438,-498436,-498434,-498432,-498431,-498429,-498427,-498425,-498423,-498421,-498420,-498418,-498416,-498414,-498412,-498410,-498408,-498407,-498405,-498403,-498401,-498399,-498397,-498395,-498394,-498392,-498390,-498388,-498386,-498384,-498382,-498381,-498379,-498377,-498375,-498373,-498371,-498370,-498368,-498366,-498364,-498362,-498360,-498358,-498357,-498355,-498353,-498351,-498349,-498347,-498345,-498344,-498342,-498340,-498338,-498336,-498334,-498332,-498331,-498329,-498327,-498325,-498323,-498321,-498319,-498318,-498316,-498314,-498312,-498310,-498308,-498306,-498305,-498303,-498301,-498299,-498297,-498295,-498293,-498292,-498290,-498288,-498286,-498284,-498282,-498280,-498279,-498277,-498275,-498273,-498271,-498269,-498267,-498265,-498264,-498262,-498260,-498258,-498256,-498254,-498252,-498251,-498249,-498247,-498245,-498243,-498241,-498239,-498238,-498236,-498234,-498232,-498230,-498228,-498226,-498225,-498223,-498221,-498219,-498217,-498215,-498213,-498211,-498210,-498208,-498206,-498204,-498202,-498200,-498198,-498197,-498195,-498193,-498191,-498189,-498187,-498185,-498183,-498182,-498180,-498178,-498176,-498174,-498172,-498170,-498169,-498167,-498165,-498163,-498161,-498159,-498157,-498155,-498154,-498152,-498150,-498148,-498146,-498144,-498142,-498140,-498139,-498137,-498135,-498133,-498131,-498129,-498127,-498126,-498124,-498122,-498120,-498118,-498116,-498114,-498112,-498111,-498109,-498107,-498105,-498103,-498101,-498099,-498097,-498096,-498094,-498092,-498090,-498088,-498086,-498084,-498082,-498081,-498079,-498077,-498075,-498073,-498071,-498069,-498067,-498066,-498064,-498062,-498060,-498058,-498056,-498054,-498052,-498051,-498049,-498047,-498045,-498043,-498041,-498039,-498037,-498036,-498034,-498032,-498030,-498028,-498026,-498024,-498022,-498021,-498019,-498017,-498015,-498013,-498011,-498009,-498007,-498005,-498004,-498002,-498000,-497998,-497996,-497994,-497992,-497990,-497989,-497987,-497985,-497983,-497981,-497979,-497977,-497975,-497974,-497972,-497970,-497968,-497966,-497964,-497962,-497960,-497958,-497957,-497955,-497953,-497951,-497949,-497947,-497945,-497943,-497942,-497940,-497938,-497936,-497934,-497932,-497930,-497928,-497926,-497925,-497923,-497921,-497919,-497917,-497915,-497913,-497911,-497909,-497908,-497906,-497904,-497902,-497900,-497898,-497896,-497894,-497892,-497891,-497889,-497887,-497885,-497883,-497881,-497879,-497877,-497875,-497874,-497872,-497870,-497868,-497866,-497864,-497862,-497860,-497858,-497857,-497855,-497853,-497851,-497849,-497847,-497845,-497843,-497841,-497840,-497838,-497836,-497834,-497832,-497830,-497828,-497826,-497824,-497823,-497821,-497819,-497817,-497815,-497813,-497811,-497809,-497807,-497805,-497804,-497802,-497800,-497798,-497796,-497794,-497792,-497790,-497788,-497787,-497785,-497783,-497781,-497779,-497777,-497775,-497773,-497771,-497769,-497768,-497766,-497764,-497762,-497760,-497758,-497756,-497754,-497752,-497751,-497749,-497747,-497745,-497743,-497741,-497739,-497737,-497735,-497733,-497732,-497730,-497728,-497726,-497724,-497722,-497720,-497718,-497716,-497714,-497713,-497711,-497709,-497707,-497705,-497703,-497701,-497699,-497697,-497695,-497694,-497692,-497690,-497688,-497686,-497684,-497682,-497680,-497678,-497676,-497675,-497673,-497671,-497669,-497667,-497665,-497663,-497661,-497659,-497657,-497655,-497654,-497652,-497650,-497648,-497646,-497644,-497642,-497640,-497638,-497636,-497635,-497633,-497631,-497629,-497627,-497625,-497623,-497621,-497619,-497617,-497615,-497614,-497612,-497610,-497608,-497606,-497604,-497602,-497600,-497598,-497596,-497594,-497593,-497591,-497589,-497587,-497585,-497583,-497581,-497579,-497577,-497575,-497573,-497572,-497570,-497568,-497566,-497564,-497562,-497560,-497558,-497556,-497554,-497552,-497551,-497549,-497547,-497545,-497543,-497541,-497539,-497537,-497535,-497533,-497531,-497529,-497528,-497526,-497524,-497522,-497520,-497518,-497516,-497514,-497512,-497510,-497508,-497507,-497505,-497503,-497501,-497499,-497497,-497495,-497493,-497491,-497489,-497487,-497485,-497484,-497482,-497480,-497478,-497476,-497474,-497472,-497470,-497468,-497466,-497464,-497462,-497461,-497459,-497457,-497455,-497453,-497451,-497449,-497447,-497445,-497443,-497441,-497439,-497437,-497436,-497434,-497432,-497430,-497428,-497426,-497424,-497422,-497420,-497418,-497416,-497414,-497413,-497411,-497409,-497407,-497405,-497403,-497401,-497399,-497397,-497395,-497393,-497391,-497389,-497388,-497386,-497384,-497382,-497380,-497378,-497376,-497374,-497372,-497370,-497368,-497366,-497364,-497363,-497361,-497359,-497357,-497355,-497353,-497351,-497349,-497347,-497345,-497343,-497341,-497339,-497337,-497336,-497334,-497332,-497330,-497328,-497326,-497324,-497322,-497320,-497318,-497316,-497314,-497312,-497311,-497309,-497307,-497305,-497303,-497301,-497299,-497297,-497295,-497293,-497291,-497289,-497287,-497285,-497284,-497282,-497280,-497278,-497276,-497274,-497272,-497270,-497268,-497266,-497264,-497262,-497260,-497258,-497256,-497255,-497253,-497251,-497249,-497247,-497245,-497243,-497241,-497239,-497237,-497235,-497233,-497231,-497229,-497227,-497226,-497224,-497222,-497220,-497218,-497216,-497214,-497212,-497210,-497208,-497206,-497204,-497202,-497200,-497198,-497197,-497195,-497193,-497191,-497189,-497187,-497185,-497183,-497181,-497179,-497177,-497175,-497173,-497171,-497169,-497167,-497166,-497164,-497162,-497160,-497158,-497156,-497154,-497152,-497150,-497148,-497146,-497144,-497142,-497140,-497138,-497136,-497134,-497133,-497131,-497129,-497127,-497125,-497123,-497121,-497119,-497117,-497115,-497113,-497111,-497109,-497107,-497105,-497103,-497101,-497100,-497098,-497096,-497094,-497092,-497090,-497088,-497086,-497084,-497082,-497080,-497078,-497076,-497074,-497072,-497070,-497068,-497066,-497065,-497063,-497061,-497059,-497057,-497055,-497053,-497051,-497049,-497047,-497045,-497043,-497041,-497039,-497037,-497035,-497033,-497031,-497029,-497028,-497026,-497024,-497022,-497020,-497018,-497016,-497014,-497012,-497010,-497008,-497006,-497004,-497002,-497000,-496998,-496996,-496994,-496992,-496991,-496989,-496987,-496985,-496983,-496981,-496979,-496977,-496975,-496973,-496971,-496969,-496967,-496965,-496963,-496961,-496959,-496957,-496955,-496953,-496951,-496950,-496948,-496946,-496944,-496942,-496940,-496938,-496936,-496934,-496932,-496930,-496928,-496926,-496924,-496922,-496920,-496918,-496916,-496914,-496912,-496910,-496908,-496907,-496905,-496903,-496901,-496899,-496897,-496895,-496893,-496891,-496889,-496887,-496885,-496883,-496881,-496879,-496877,-496875,-496873,-496871,-496869,-496867,-496865,-496863,-496862,-496860,-496858,-496856,-496854,-496852,-496850,-496848,-496846,-496844,-496842,-496840,-496838,-496836,-496834,-496832,-496830,-496828,-496826,-496824,-496822,-496820,-496818,-496816,-496814,-496812,-496811,-496809,-496807,-496805,-496803,-496801,-496799,-496797,-496795,-496793,-496791,-496789,-496787,-496785,-496783,-496781,-496779,-496777,-496775,-496773,-496771,-496769,-496767,-496765,-496763,-496761,-496759,-496757,-496756,-496754,-496752,-496750,-496748,-496746,-496744,-496742,-496740,-496738,-496736,-496734,-496732,-496730,-496728,-496726,-496724,-496722,-496720,-496718,-496716,-496714,-496712,-496710,-496708,-496706,-496704,-496702,-496700,-496698,-496696,-496694,-496693,-496691,-496689,-496687,-496685,-496683,-496681,-496679,-496677,-496675,-496673,-496671,-496669,-496667,-496665,-496663,-496661,-496659,-496657,-496655,-496653,-496651,-496649,-496647,-496645,-496643,-496641,-496639,-496637,-496635,-496633,-496631,-496629,-496627,-496625,-496623,-496621,-496620,-496618,-496616,-496614,-496612,-496610,-496608,-496606,-496604,-496602,-496600,-496598,-496596,-496594,-496592,-496590,-496588,-496586,-496584,-496582,-496580,-496578,-496576,-496574,-496572,-496570,-496568,-496566,-496564,-496562,-496560,-496558,-496556,-496554,-496552,-496550,-496548,-496546,-496544,-496542,-496540,-496538,-496536,-496534,-496532,-496530,-496529,-496527,-496525,-496523,-496521,-496519,-496517,-496515,-496513,-496511,-496509,-496507,-496505,-496503,-496501,-496499,-496497,-496495,-496493,-496491,-496489,-496487,-496485,-496483,-496481,-496479,-496477,-496475,-496473,-496471,-496469,-496467,-496465,-496463,-496461,-496459,-496457,-496455,-496453,-496451,-496449,-496447,-496445,-496443,-496441,-496439,-496437,-496435,-496433,-496431,-496429,-496427,-496425,-496423,-496421,-496419,-496417,-496415,-496413,-496411,-496409,-496407,-496405,-496403,-496401,-496399,-496397,-496395,-496393,-496391,-496389,-496387,-496385,-496383,-496382,-496380,-496378,-496376,-496374,-496372,-496370,-496368,-496366,-496364,-496362,-496360,-496358,-496356,-496354,-496352,-496350,-496348,-496346,-496344,-496342,-496340,-496338,-496336,-496334,-496332,-496330,-496328,-496326,-496324,-496322,-496320,-496318,-496316,-496314,-496312,-496310,-496308,-496306,-496304,-496302,-496300,-496298,-496296,-496294,-496292,-496290,-496288,-496286,-496284,-496282,-496280,-496278,-496276,-496274,-496272,-496270,-496268,-496266,-496264,-496262,-496260,-496258,-496256,-496254,-496252,-496250,-496248,-496246,-496244,-496242,-496240,-496238,-496236,-496234,-496232,-496230,-496228,-496226,-496224,-496222,-496220,-496218,-496216,-496214,-496212,-496210,-496208,-496206,-496204,-496202,-496200,-496198,-496196,-496194,-496192,-496190,-496188,-496186,-496184,-496182,-496180,-496178,-496176,-496174,-496172,-496170,-496168,-496166,-496164,-496162,-496160,-496158,-496156,-496154,-496152,-496150,-496148,-496146,-496144,-496142,-496140,-496138,-496136,-496134,-496132,-496130,-496128,-496126,-496124,-496121,-496119,-496117,-496115,-496113,-496111,-496109,-496107,-496105,-496103,-496101,-496099,-496097,-496095,-496093,-496091,-496089,-496087,-496085,-496083,-496081,-496079,-496077,-496075,-496073,-496071,-496069,-496067,-496065,-496063,-496061,-496059,-496057,-496055,-496053,-496051,-496049,-496047,-496045,-496043,-496041,-496039,-496037,-496035,-496033,-496031,-496029,-496027,-496025,-496023,-496021,-496019,-496017,-496015,-496013,-496011,-496009,-496007,-496005,-496003,-496001,-495999,-495997,-495995,-495993,-495991,-495989,-495987,-495985,-495983,-495981,-495979,-495977,-495975,-495972,-495970,-495968,-495966,-495964,-495962,-495960,-495958,-495956,-495954,-495952,-495950,-495948,-495946,-495944,-495942,-495940,-495938,-495936,-495934,-495932,-495930,-495928,-495926,-495924,-495922,-495920,-495918,-495916,-495914,-495912,-495910,-495908,-495906,-495904,-495902,-495900,-495898,-495896,-495894,-495892,-495890,-495888,-495886,-495884,-495882,-495879,-495877,-495875,-495873,-495871,-495869,-495867,-495865,-495863,-495861,-495859,-495857,-495855,-495853,-495851,-495849,-495847,-495845,-495843,-495841,-495839,-495837,-495835,-495833,-495831,-495829,-495827,-495825,-495823,-495821,-495819,-495817,-495815,-495813,-495811,-495809,-495807,-495804,-495802,-495800,-495798,-495796,-495794,-495792,-495790,-495788,-495786,-495784,-495782,-495780,-495778,-495776,-495774,-495772,-495770,-495768,-495766,-495764,-495762,-495760,-495758,-495756,-495754,-495752,-495750,-495748,-495746,-495744,-495742,-495739,-495737,-495735,-495733,-495731,-495729,-495727,-495725,-495723,-495721,-495719,-495717,-495715,-495713,-495711,-495709,-495707,-495705,-495703,-495701,-495699,-495697,-495695,-495693,-495691,-495689,-495687,-495685,-495682,-495680,-495678,-495676,-495674,-495672,-495670,-495668,-495666,-495664,-495662,-495660,-495658,-495656,-495654,-495652,-495650,-495648,-495646,-495644,-495642,-495640,-495638,-495636,-495634,-495632,-495629,-495627,-495625,-495623,-495621,-495619,-495617,-495615,-495613,-495611,-495609,-495607,-495605,-495603,-495601,-495599,-495597,-495595,-495593,-495591,-495589,-495587,-495585,-495582,-495580,-495578,-495576,-495574,-495572,-495570,-495568,-495566,-495564,-495562,-495560,-495558,-495556,-495554,-495552,-495550,-495548,-495546,-495544,-495542,-495540,-495537,-495535,-495533,-495531,-495529,-495527,-495525,-495523,-495521,-495519,-495517,-495515,-495513,-495511,-495509,-495507,-495505,-495503,-495501,-495499,-495497,-495494,-495492,-495490,-495488,-495486,-495484,-495482,-495480,-495478,-495476,-495474,-495472,-495470,-495468,-495466,-495464,-495462,-495460,-495458,-495456,-495453,-495451,-495449,-495447,-495445,-495443,-495441,-495439,-495437,-495435,-495433,-495431,-495429,-495427,-495425,-495423,-495421,-495419,-495416,-495414,-495412,-495410,-495408,-495406,-495404,-495402,-495400,-495398,-495396,-495394,-495392,-495390,-495388,-495386,-495384,-495382,-495379,-495377,-495375,-495373,-495371,-495369,-495367,-495365,-495363,-495361,-495359,-495357,-495355,-495353,-495351,-495349,-495347,-495344,-495342,-495340,-495338,-495336,-495334,-495332,-495330,-495328,-495326,-495324,-495322,-495320,-495318,-495316,-495314,-495312,-495309,-495307,-495305,-495303,-495301,-495299,-495297,-495295,-495293,-495291,-495289,-495287,-495285,-495283,-495281,-495279,-495276,-495274,-495272,-495270,-495268,-495266,-495264,-495262,-495260,-495258,-495256,-495254,-495252,-495250,-495248,-495245,-495243,-495241,-495239,-495237,-495235,-495233,-495231,-495229,-495227,-495225,-495223,-495221,-495219,-495217,-495214,-495212,-495210,-495208,-495206,-495204,-495202,-495200,-495198,-495196,-495194,-495192,-495190,-495188,-495186,-495183,-495181,-495179,-495177,-495175,-495173,-495171,-495169,-495167,-495165,-495163,-495161,-495159,-495157,-495154,-495152,-495150,-495148,-495146,-495144,-495142,-495140,-495138,-495136,-495134,-495132,-495130,-495128,-495125,-495123,-495121,-495119,-495117,-495115,-495113,-495111,-495109,-495107,-495105,-495103,-495101,-495098,-495096,-495094,-495092,-495090,-495088,-495086,-495084,-495082,-495080,-495078,-495076,-495074,-495071,-495069,-495067,-495065,-495063,-495061,-495059,-495057,-495055,-495053,-495051,-495049,-495047,-495044,-495042,-495040,-495038,-495036,-495034,-495032,-495030,-495028,-495026,-495024,-495022,-495020,-495017,-495015,-495013,-495011,-495009,-495007,-495005,-495003,-495001,-494999,-494997,-494995,-494992,-494990,-494988,-494986,-494984,-494982,-494980,-494978,-494976,-494974,-494972,-494970,-494967,-494965,-494963,-494961,-494959,-494957,-494955,-494953,-494951,-494949,-494947,-494945,-494942,-494940,-494938,-494936,-494934,-494932,-494930,-494928,-494926,-494924,-494922,-494920,-494917,-494915,-494913,-494911,-494909,-494907,-494905,-494903,-494901,-494899,-494897,-494894,-494892,-494890,-494888,-494886,-494884,-494882,-494880,-494878,-494876,-494874,-494871,-494869,-494867,-494865,-494863,-494861,-494859,-494857,-494855,-494853,-494851,-494849,-494846,-494844,-494842,-494840,-494838,-494836,-494834,-494832,-494830,-494828,-494825,-494823,-494821,-494819,-494817,-494815,-494813,-494811,-494809,-494807,-494805,-494802,-494800,-494798,-494796,-494794,-494792,-494790,-494788,-494786,-494784,-494782,-494779,-494777,-494775,-494773,-494771,-494769,-494767,-494765,-494763,-494761,-494758,-494756,-494754,-494752,-494750,-494748,-494746,-494744,-494742,-494740,-494737,-494735,-494733,-494731,-494729,-494727,-494725,-494723,-494721,-494719,-494716,-494714,-494712,-494710,-494708,-494706,-494704,-494702,-494700,-494698,-494695,-494693,-494691,-494689,-494687,-494685,-494683,-494681,-494679,-494677,-494674,-494672,-494670,-494668,-494666,-494664,-494662,-494660,-494658,-494656,-494653,-494651,-494649,-494647,-494645,-494643,-494641,-494639,-494637,-494635,-494632,-494630,-494628,-494626,-494624,-494622,-494620,-494618,-494616,-494613,-494611,-494609,-494607,-494605,-494603,-494601,-494599,-494597,-494595,-494592,-494590,-494588,-494586,-494584,-494582,-494580,-494578,-494576,-494573,-494571,-494569,-494567,-494565,-494563,-494561,-494559,-494557,-494554,-494552,-494550,-494548,-494546,-494544,-494542,-494540,-494538,-494535,-494533,-494531,-494529,-494527,-494525,-494523,-494521,-494519,-494516,-494514,-494512,-494510,-494508,-494506,-494504,-494502,-494500,-494497,-494495,-494493,-494491,-494489,-494487,-494485,-494483,-494481,-494478,-494476,-494474,-494472,-494470,-494468,-494466,-494464,-494461,-494459,-494457,-494455,-494453,-494451,-494449,-494447,-494445,-494442,-494440,-494438,-494436,-494434,-494432,-494430,-494428,-494426,-494423,-494421,-494419,-494417,-494415,-494413,-494411,-494409,-494406,-494404,-494402,-494400,-494398,-494396,-494394,-494392,-494389,-494387,-494385,-494383,-494381,-494379,-494377,-494375,-494373,-494370,-494368,-494366,-494364,-494362,-494360,-494358,-494356,-494353,-494351,-494349,-494347,-494345,-494343,-494341,-494339,-494336,-494334,-494332,-494330,-494328,-494326,-494324,-494322,-494319,-494317,-494315,-494313,-494311,-494309,-494307,-494305,-494302,-494300,-494298,-494296,-494294,-494292,-494290,-494288,-494285,-494283,-494281,-494279,-494277,-494275,-494273,-494271,-494268,-494266,-494264,-494262,-494260,-494258,-494256,-494254,-494251,-494249,-494247,-494245,-494243,-494241,-494239,-494237,-494234,-494232,-494230,-494228,-494226,-494224,-494222,-494219,-494217,-494215,-494213,-494211,-494209,-494207,-494205,-494202,-494200,-494198,-494196,-494194,-494192,-494190,-494188,-494185,-494183,-494181,-494179,-494177,-494175,-494173,-494170,-494168,-494166,-494164,-494162,-494160,-494158,-494155,-494153,-494151,-494149,-494147,-494145,-494143,-494141,-494138,-494136,-494134,-494132,-494130,-494128,-494126,-494123,-494121,-494119,-494117,-494115,-494113,-494111,-494109,-494106,-494104,-494102,-494100,-494098,-494096,-494094,-494091,-494089,-494087,-494085,-494083,-494081,-494079,-494076,-494074,-494072,-494070,-494068,-494066,-494064,-494061,-494059,-494057,-494055,-494053,-494051,-494049,-494046,-494044,-494042,-494040,-494038,-494036,-494034,-494031,-494029,-494027,-494025,-494023,-494021,-494019,-494016,-494014,-494012,-494010,-494008,-494006,-494004,-494001,-493999,-493997,-493995,-493993,-493991,-493989,-493986,-493984,-493982,-493980,-493978,-493976,-493974,-493971,-493969,-493967,-493965,-493963,-493961,-493959,-493956,-493954,-493952,-493950,-493948,-493946,-493944,-493941,-493939,-493937,-493935,-493933,-493931,-493928,-493926,-493924,-493922,-493920,-493918,-493916,-493913,-493911,-493909,-493907,-493905,-493903,-493901,-493898,-493896,-493894,-493892,-493890,-493888,-493886,-493883,-493881,-493879,-493877,-493875,-493873,-493870,-493868,-493866,-493864,-493862,-493860,-493858,-493855,-493853,-493851,-493849,-493847,-493845,-493842,-493840,-493838,-493836,-493834,-493832,-493830,-493827,-493825,-493823,-493821,-493819,-493817,-493814,-493812,-493810,-493808,-493806,-493804,-493802,-493799,-493797,-493795,-493793,-493791,-493789,-493786,-493784,-493782,-493780,-493778,-493776,-493773,-493771,-493769,-493767,-493765,-493763,-493761,-493758,-493756,-493754,-493752,-493750,-493748,-493745,-493743,-493741,-493739,-493737,-493735,-493732,-493730,-493728,-493726,-493724,-493722,-493719,-493717,-493715,-493713,-493711,-493709,-493706,-493704,-493702,-493700,-493698,-493696,-493694,-493691,-493689,-493687,-493685,-493683,-493681,-493678,-493676,-493674,-493672,-493670,-493668,-493665,-493663,-493661,-493659,-493657,-493655,-493652,-493650,-493648,-493646,-493644,-493642,-493639,-493637,-493635,-493633,-493631,-493629,-493626,-493624,-493622,-493620,-493618,-493616,-493613,-493611,-493609,-493607,-493605,-493603,-493600,-493598,-493596,-493594,-493592,-493590,-493587,-493585,-493583,-493581,-493579,-493577,-493574,-493572,-493570,-493568,-493566,-493564,-493561,-493559,-493557,-493555,-493553,-493550,-493548,-493546,-493544,-493542,-493540,-493537,-493535,-493533,-493531,-493529,-493527,-493524,-493522,-493520,-493518,-493516,-493514,-493511,-493509,-493507,-493505,-493503,-493500,-493498,-493496,-493494,-493492,-493490,-493487,-493485,-493483,-493481,-493479,-493477,-493474,-493472,-493470,-493468,-493466,-493464,-493461,-493459,-493457,-493455,-493453,-493450,-493448,-493446,-493444,-493442,-493440,-493437,-493435,-493433,-493431,-493429,-493426,-493424,-493422,-493420,-493418,-493416,-493413,-493411,-493409,-493407,-493405,-493403,-493400,-493398,-493396,-493394,-493392,-493389,-493387,-493385,-493383,-493381,-493379,-493376,-493374,-493372,-493370,-493368,-493365,-493363,-493361,-493359,-493357,-493354,-493352,-493350,-493348,-493346,-493344,-493341,-493339,-493337,-493335,-493333,-493330,-493328,-493326,-493324,-493322,-493320,-493317,-493315,-493313,-493311,-493309,-493306,-493304,-493302,-493300,-493298,-493295,-493293,-493291,-493289,-493287,-493285,-493282,-493280,-493278,-493276,-493274,-493271,-493269,-493267,-493265,-493263,-493260,-493258,-493256,-493254,-493252,-493250,-493247,-493245,-493243,-493241,-493239,-493236,-493234,-493232,-493230,-493228,-493225,-493223,-493221,-493219,-493217,-493214,-493212,-493210,-493208,-493206,-493204,-493201,-493199,-493197,-493195,-493193,-493190,-493188,-493186,-493184,-493182,-493179,-493177,-493175,-493173,-493171,-493168,-493166,-493164,-493162,-493160,-493157,-493155,-493153,-493151,-493149,-493146,-493144,-493142,-493140,-493138,-493135,-493133,-493131,-493129,-493127,-493124,-493122,-493120,-493118,-493116,-493114,-493111,-493109,-493107,-493105,-493103,-493100,-493098,-493096,-493094,-493092,-493089,-493087,-493085,-493083,-493081,-493078,-493076,-493074,-493072,-493070,-493067,-493065,-493063,-493061,-493059,-493056,-493054,-493052,-493050,-493048,-493045,-493043,-493041,-493039,-493036,-493034,-493032,-493030,-493028,-493025,-493023,-493021,-493019,-493017,-493014,-493012,-493010,-493008,-493006,-493003,-493001,-492999,-492997,-492995,-492992,-492990,-492988,-492986,-492984,-492981,-492979,-492977,-492975,-492973,-492970,-492968,-492966,-492964,-492962,-492959,-492957,-492955,-492953,-492950,-492948,-492946,-492944,-492942,-492939,-492937,-492935,-492933,-492931,-492928,-492926,-492924,-492922,-492920,-492917,-492915,-492913,-492911,-492909,-492906,-492904,-492902,-492900,-492897,-492895,-492893,-492891,-492889,-492886,-492884,-492882,-492880,-492878,-492875,-492873,-492871,-492869,-492866,-492864,-492862,-492860,-492858,-492855,-492853,-492851,-492849,-492847,-492844,-492842,-492840,-492838,-492835,-492833,-492831,-492829,-492827,-492824,-492822,-492820,-492818,-492816,-492813,-492811,-492809,-492807,-492804,-492802,-492800,-492798,-492796,-492793,-492791,-492789,-492787,-492785,-492782,-492780,-492778,-492776,-492773,-492771,-492769,-492767,-492765,-492762,-492760,-492758,-492756,-492753,-492751,-492749,-492747,-492745,-492742,-492740,-492738,-492736,-492733,-492731,-492729,-492727,-492725,-492722,-492720,-492718,-492716,-492713,-492711,-492709,-492707,-492705,-492702,-492700,-492698,-492696,-492693,-492691,-492689,-492687,-492685,-492682,-492680,-492678,-492676,-492673,-492671,-492669,-492667,-492665,-492662,-492660,-492658,-492656,-492653,-492651,-492649,-492647,-492645,-492642,-492640,-492638,-492636,-492633,-492631,-492629,-492627,-492625,-492622,-492620,-492618,-492616,-492613,-492611,-492609,-492607,-492604,-492602,-492600,-492598,-492596,-492593,-492591,-492589,-492587,-492584,-492582,-492580,-492578,-492575,-492573,-492571,-492569,-492567,-492564,-492562,-492560,-492558,-492555,-492553,-492551,-492549,-492546,-492544,-492542,-492540,-492538,-492535,-492533,-492531,-492529,-492526,-492524,-492522,-492520,-492517,-492515,-492513,-492511,-492509,-492506,-492504,-492502,-492500,-492497,-492495,-492493,-492491,-492488,-492486,-492484,-492482,-492479,-492477,-492475,-492473,-492471,-492468,-492466,-492464,-492462,-492459,-492457,-492455,-492453,-492450,-492448,-492446,-492444,-492441,-492439,-492437,-492435,-492432,-492430,-492428,-492426,-492424,-492421,-492419,-492417,-492415,-492412,-492410,-492408,-492406,-492403,-492401,-492399,-492397,-492394,-492392,-492390,-492388,-492385,-492383,-492381,-492379,-492376,-492374,-492372,-492370,-492367,-492365,-492363,-492361,-492359,-492356,-492354,-492352,-492350,-492347,-492345,-492343,-492341,-492338,-492336,-492334,-492332,-492329,-492327,-492325,-492323,-492320,-492318,-492316,-492314,-492311,-492309,-492307,-492305,-492302,-492300,-492298,-492296,-492293,-492291,-492289,-492287,-492284,-492282,-492280,-492278,-492275,-492273,-492271,-492269,-492266,-492264,-492262,-492260,-492257,-492255,-492253,-492251,-492248,-492246,-492244,-492242,-492239,-492237,-492235,-492233,-492230,-492228,-492226,-492224,-492221,-492219,-492217,-492215,-492212,-492210,-492208,-492206,-492203,-492201,-492199,-492197,-492194,-492192,-492190,-492188,-492185,-492183,-492181,-492179,-492176,-492174,-492172,-492170,-492167,-492165,-492163,-492161,-492158,-492156,-492154,-492152,-492149,-492147,-492145,-492143,-492140,-492138,-492136,-492134,-492131,-492129,-492127,-492125,-492122,-492120,-492118,-492116,-492113,-492111,-492109,-492106,-492104,-492102,-492100,-492097,-492095,-492093,-492091,-492088,-492086,-492084,-492082,-492079,-492077,-492075,-492073,-492070,-492068,-492066,-492064,-492061,-492059,-492057,-492055,-492052,-492050,-492048,-492045,-492043,-492041,-492039,-492036,-492034,-492032,-492030,-492027,-492025,-492023,-492021,-492018,-492016,-492014,-492012,-492009,-492007,-492005,-492002,-492000,-491998,-491996,-491993,-491991,-491989,-491987,-491984,-491982,-491980,-491978,-491975,-491973,-491971,-491969,-491966,-491964,-491962,-491959,-491957,-491955,-491953,-491950,-491948,-491946,-491944,-491941,-491939,-491937,-491935,-491932,-491930,-491928,-491925,-491923,-491921,-491919,-491916,-491914,-491912,-491910,-491907,-491905,-491903,-491900,-491898,-491896,-491894,-491891,-491889,-491887,-491885,-491882,-491880,-491878,-491876,-491873,-491871,-491869,-491866,-491864,-491862,-491860,-491857,-491855,-491853,-491851,-491848,-491846,-491844,-491841,-491839,-491837,-491835,-491832,-491830,-491828,-491826,-491823,-491821,-491819,-491816,-491814,-491812,-491810,-491807,-491805,-491803,-491801,-491798,-491796,-491794,-491791,-491789,-491787,-491785,-491782,-491780,-491778,-491775,-491773,-491771,-491769,-491766,-491764,-491762,-491760,-491757,-491755,-491753,-491750,-491748,-491746,-491744,-491741,-491739,-491737,-491734,-491732,-491730,-491728,-491725,-491723,-491721,-491718,-491716,-491714,-491712,-491709,-491707,-491705,-491703,-491700,-491698,-491696,-491693,-491691,-491689,-491687,-491684,-491682,-491680,-491677,-491675,-491673,-491671,-491668,-491666,-491664,-491661,-491659,-491657,-491655,-491652,-491650,-491648,-491645,-491643,-491641,-491639,-491636,-491634,-491632,-491629,-491627,-491625,-491623,-491620,-491618,-491616,-491613,-491611,-491609,-491607,-491604,-491602,-491600,-491597,-491595,-491593,-491591,-491588,-491586,-491584,-491581,-491579,-491577,-491575,-491572,-491570,-491568,-491565,-491563,-491561,-491559,-491556,-491554,-491552,-491549,-491547,-491545,-491543,-491540,-491538,-491536,-491533,-491531,-491529,-491526,-491524,-491522,-491520,-491517,-491515,-491513,-491510,-491508,-491506,-491504,-491501,-491499,-491497,-491494,-491492,-491490,-491488,-491485,-491483,-491481,-491478,-491476,-491474,-491471,-491469,-491467,-491465,-491462,-491460,-491458,-491455,-491453,-491451,-491449,-491446,-491444,-491442,-491439,-491437,-491435,-491432,-491430,-491428,-491426,-491423,-491421,-491419,-491416,-491414,-491412,-491409,-491407,-491405,-491403,-491400,-491398,-491396,-491393,-491391,-491389,-491386,-491384,-491382,-491380,-491377,-491375,-491373,-491370,-491368,-491366,-491363,-491361,-491359,-491357,-491354,-491352,-491350,-491347,-491345,-491343,-491340,-491338,-491336,-491334,-491331,-491329,-491327,-491324,-491322,-491320,-491317,-491315,-491313,-491311,-491308,-491306,-491304,-491301,-491299,-491297,-491294,-491292,-491290,-491287,-491285,-491283,-491281,-491278,-491276,-491274,-491271,-491269,-491267,-491264,-491262,-491260,-491258,-491255,-491253,-491251,-491248,-491246,-491244,-491241,-491239,-491237,-491234,-491232,-491230,-491228,-491225,-491223,-491221,-491218,-491216,-491214,-491211,-491209,-491207,-491204,-491202,-491200,-491197,-491195,-491193,-491191,-491188,-491186,-491184,-491181,-491179,-491177,-491174,-491172,-491170,-491167,-491165,-491163,-491161,-491158,-491156,-491154,-491151,-491149,-491147,-491144,-491142,-491140,-491137,-491135,-491133,-491130,-491128,-491126,-491124,-491121,-491119,-491117,-491114,-491112,-491110,-491107,-491105,-491103,-491100,-491098,-491096,-491093,-491091,-491089,-491086,-491084,-491082,-491080,-491077,-491075,-491073,-491070,-491068,-491066,-491063,-491061,-491059,-491056,-491054,-491052,-491049,-491047,-491045,-491042,-491040,-491038,-491035,-491033,-491031,-491029,-491026,-491024,-491022,-491019,-491017,-491015,-491012,-491010,-491008,-491005,-491003,-491001,-490998,-490996,-490994,-490991,-490989,-490987,-490984,-490982,-490980,-490977,-490975,-490973,-490970,-490968,-490966,-490964,-490961,-490959,-490957,-490954,-490952,-490950,-490947,-490945,-490943,-490940,-490938,-490936,-490933,-490931,-490929,-490926,-490924,-490922,-490919,-490917,-490915,-490912,-490910,-490908,-490905,-490903,-490901,-490898,-490896,-490894,-490891,-490889,-490887,-490884,-490882,-490880,-490877,-490875,-490873,-490870,-490868,-490866,-490863,-490861,-490859,-490856,-490854,-490852,-490850,-490847,-490845,-490843,-490840,-490838,-490836,-490833,-490831,-490829,-490826,-490824,-490822,-490819,-490817,-490815,-490812,-490810,-490808,-490805,-490803,-490801,-490798,-490796,-490794,-490791,-490789,-490787,-490784,-490782,-490780,-490777,-490775,-490773,-490770,-490768,-490766,-490763,-490761,-490759,-490756,-490754,-490752,-490749,-490747,-490745,-490742,-490740,-490738,-490735,-490733,-490731,-490728,-490726,-490724,-490721,-490719,-490716,-490714,-490712,-490709,-490707,-490705,-490702,-490700,-490698,-490695,-490693,-490691,-490688,-490686,-490684,-490681,-490679,-490677,-490674,-490672,-490670,-490667,-490665,-490663,-490660,-490658,-490656,-490653,-490651,-490649,-490646,-490644,-490642,-490639,-490637,-490635,-490632,-490630,-490628,-490625,-490623,-490621,-490618,-490616,-490614,-490611,-490609,-490606,-490604,-490602,-490599,-490597,-490595,-490592,-490590,-490588,-490585,-490583,-490581,-490578,-490576,-490574,-490571,-490569,-490567,-490564,-490562,-490560,-490557,-490555,-490553,-490550,-490548,-490546,-490543,-490541,-490538,-490536,-490534,-490531,-490529,-490527,-490524,-490522,-490520,-490517,-490515,-490513,-490510,-490508,-490506,-490503,-490501,-490499,-490496,-490494,-490492,-490489,-490487,-490484,-490482,-490480,-490477,-490475,-490473,-490470,-490468,-490466,-490463,-490461,-490459,-490456,-490454,-490452,-490449,-490447,-490444,-490442,-490440,-490437,-490435,-490433,-490430,-490428,-490426,-490423,-490421,-490419,-490416,-490414,-490412,-490409,-490407,-490404,-490402,-490400,-490397,-490395,-490393,-490390,-490388,-490386,-490383,-490381,-490379,-490376,-490374,-490371,-490369,-490367,-490364,-490362,-490360,-490357,-490355,-490353,-490350,-490348,-490346,-490343,-490341,-490338,-490336,-490334,-490331,-490329,-490327,-490324,-490322,-490320,-490317,-490315,-490313,-490310,-490308,-490305,-490303,-490301,-490298,-490296,-490294,-490291,-490289,-490287,-490284,-490282,-490279,-490277,-490275,-490272,-490270,-490268,-490265,-490263,-490261,-490258,-490256,-490253,-490251,-490249,-490246,-490244,-490242,-490239,-490237,-490235,-490232,-490230,-490227,-490225,-490223,-490220,-490218,-490216,-490213,-490211,-490209,-490206,-490204,-490201,-490199,-490197,-490194,-490192,-490190,-490187,-490185,-490183,-490180,-490178,-490175,-490173,-490171,-490168,-490166,-490164,-490161,-490159,-490156,-490154,-490152,-490149,-490147,-490145,-490142,-490140,-490138,-490135,-490133,-490130,-490128,-490126,-490123,-490121,-490119,-490116,-490114,-490111,-490109,-490107,-490104,-490102,-490100,-490097,-490095,-490093,-490090,-490088,-490085,-490083,-490081,-490078,-490076,-490074,-490071,-490069,-490066,-490064,-490062,-490059,-490057,-490055,-490052,-490050,-490047,-490045,-490043,-490040,-490038,-490036,-490033,-490031,-490028,-490026,-490024,-490021,-490019,-490017,-490014,-490012,-490009,-490007,-490005,-490002,-490000,-489998,-489995,-489993,-489990,-489988,-489986,-489983,-489981,-489978,-489976,-489974,-489971,-489969,-489967,-489964,-489962,-489959,-489957,-489955,-489952,-489950,-489948,-489945,-489943,-489940,-489938,-489936,-489933,-489931,-489929,-489926,-489924,-489921,-489919,-489917,-489914,-489912,-489909,-489907,-489905,-489902,-489900,-489898,-489895,-489893,-489890,-489888,-489886,-489883,-489881,-489878,-489876,-489874,-489871,-489869,-489867,-489864,-489862,-489859,-489857,-489855,-489852,-489850,-489847,-489845,-489843,-489840,-489838,-489836,-489833,-489831,-489828,-489826,-489824,-489821,-489819,-489816,-489814,-489812,-489809,-489807,-489805,-489802,-489800,-489797,-489795,-489793,-489790,-489788,-489785,-489783,-489781,-489778,-489776,-489773,-489771,-489769,-489766,-489764,-489762,-489759,-489757,-489754,-489752,-489750,-489747,-489745,-489742,-489740,-489738,-489735,-489733,-489730,-489728,-489726,-489723,-489721,-489718,-489716,-489714,-489711,-489709,-489707,-489704,-489702,-489699,-489697,-489695,-489692,-489690,-489687,-489685,-489683,-489680,-489678,-489675,-489673,-489671,-489668,-489666,-489663,-489661,-489659,-489656,-489654,-489651,-489649,-489647,-489644,-489642,-489639,-489637,-489635,-489632,-489630,-489627,-489625,-489623,-489620,-489618,-489615,-489613,-489611,-489608,-489606,-489603,-489601,-489599,-489596,-489594,-489591,-489589,-489587,-489584,-489582,-489579,-489577,-489575,-489572,-489570,-489567,-489565,-489563,-489560,-489558,-489555,-489553,-489551,-489548,-489546,-489543,-489541,-489539,-489536,-489534,-489531,-489529,-489527,-489524,-489522,-489519,-489517,-489515,-489512,-489510,-489507,-489505,-489503,-489500,-489498,-489495,-489493,-489491,-489488,-489486,-489483,-489481,-489479,-489476,-489474,-489471,-489469,-489467,-489464,-489462,-489459,-489457,-489454,-489452,-489450,-489447,-489445,-489442,-489440,-489438,-489435,-489433,-489430,-489428,-489426,-489423,-489421,-489418,-489416,-489414,-489411,-489409,-489406,-489404,-489401,-489399,-489397,-489394,-489392,-489389,-489387,-489385,-489382,-489380,-489377,-489375,-489373,-489370,-489368,-489365,-489363,-489361,-489358,-489356,-489353,-489351,-489348,-489346,-489344,-489341,-489339,-489336,-489334,-489332,-489329,-489327,-489324,-489322,-489319,-489317,-489315,-489312,-489310,-489307,-489305,-489303,-489300,-489298,-489295,-489293,-489290,-489288,-489286,-489283,-489281,-489278,-489276,-489274,-489271,-489269,-489266,-489264,-489261,-489259,-489257,-489254,-489252,-489249,-489247,-489245,-489242,-489240,-489237,-489235,-489232,-489230,-489228,-489225,-489223,-489220,-489218,-489216,-489213,-489211,-489208,-489206,-489203,-489201,-489199,-489196,-489194,-489191,-489189,-489186,-489184,-489182,-489179,-489177,-489174,-489172,-489170,-489167,-489165,-489162,-489160,-489157,-489155,-489153,-489150,-489148,-489145,-489143,-489140,-489138,-489136,-489133,-489131,-489128,-489126,-489123,-489121,-489119,-489116,-489114,-489111,-489109,-489106,-489104,-489102,-489099,-489097,-489094,-489092,-489090,-489087,-489085,-489082,-489080,-489077,-489075,-489073,-489070,-489068,-489065,-489063,-489060,-489058,-489056,-489053,-489051,-489048,-489046,-489043,-489041,-489039,-489036,-489034,-489031,-489029,-489026,-489024,-489022,-489019,-489017,-489014,-489012,-489009,-489007,-489004,-489002,-489000,-488997,-488995,-488992,-488990,-488987,-488985,-488983,-488980,-488978,-488975,-488973,-488970,-488968,-488966,-488963,-488961,-488958,-488956,-488953,-488951,-488949,-488946,-488944,-488941,-488939,-488936,-488934,-488931,-488929,-488927,-488924,-488922,-488919,-488917,-488914,-488912,-488910,-488907,-488905,-488902,-488900,-488897,-488895,-488893,-488890,-488888,-488885,-488883,-488880,-488878,-488875,-488873,-488871,-488868,-488866,-488863,-488861,-488858,-488856,-488853,-488851,-488849,-488846,-488844,-488841,-488839,-488836,-488834,-488832,-488829,-488827,-488824,-488822,-488819,-488817,-488814,-488812,-488810,-488807,-488805,-488802,-488800,-488797,-488795,-488792,-488790,-488788,-488785,-488783,-488780,-488778,-488775,-488773,-488770,-488768,-488766,-488763,-488761,-488758,-488756,-488753,-488751,-488748,-488746,-488744,-488741,-488739,-488736,-488734,-488731,-488729,-488726,-488724,-488722,-488719,-488717,-488714,-488712,-488709,-488707,-488704,-488702,-488700,-488697,-488695,-488692,-488690,-488687,-488685,-488682,-488680,-488678,-488675,-488673,-488670,-488668,-488665,-488663,-488660,-488658,-488655,-488653,-488651,-488648,-488646,-488643,-488641,-488638,-488636,-488633,-488631,-488628,-488626,-488624,-488621,-488619,-488616,-488614,-488611,-488609,-488606,-488604,-488602,-488599,-488597,-488594,-488592,-488589,-488587,-488584,-488582,-488579,-488577,-488575,-488572,-488570,-488567,-488565,-488562,-488560,-488557,-488555,-488552,-488550,-488548,-488545,-488543,-488540,-488538,-488535,-488533,-488530,-488528,-488525,-488523,-488520,-488518,-488516,-488513,-488511,-488508,-488506,-488503,-488501,-488498,-488496,-488493,-488491,-488489,-488486,-488484,-488481,-488479,-488476,-488474,-488471,-488469,-488466,-488464,-488461,-488459,-488457,-488454,-488452,-488449,-488447,-488444,-488442,-488439,-488437,-488434,-488432,-488429,-488427,-488425,-488422,-488420,-488417,-488415,-488412,-488410,-488407,-488405,-488402,-488400,-488397,-488395,-488393,-488390,-488388,-488385,-488383,-488380,-488378,-488375,-488373,-488370,-488368,-488365,-488363,-488360,-488358,-488356,-488353,-488351,-488348,-488346,-488343,-488341,-488338,-488336,-488333,-488331,-488328,-488326,-488323,-488321,-488319,-488316,-488314,-488311,-488309,-488306,-488304,-488301,-488299,-488296,-488294,-488291,-488289,-488286,-488284,-488282,-488279,-488277,-488274,-488272,-488269,-488267,-488264,-488262,-488259,-488257,-488254,-488252,-488249,-488247,-488244,-488242,-488240,-488237,-488235,-488232,-488230,-488227,-488225,-488222,-488220,-488217,-488215,-488212,-488210,-488207,-488205,-488202,-488200,-488197,-488195,-488193,-488190,-488188,-488185,-488183,-488180,-488178,-488175,-488173,-488170,-488168,-488165,-488163,-488160,-488158,-488155,-488153,-488150,-488148,-488145,-488143,-488141,-488138,-488136,-488133,-488131,-488128,-488126,-488123,-488121,-488118,-488116,-488113,-488111,-488108,-488106,-488103,-488101,-488098,-488096,-488093,-488091,-488088,-488086,-488083,-488081,-488079,-488076,-488074,-488071,-488069,-488066,-488064,-488061,-488059,-488056,-488054,-488051,-488049,-488046,-488044,-488041,-488039,-488036,-488034,-488031,-488029,-488026,-488024,-488021,-488019,-488016,-488014,-488012,-488009,-488007,-488004,-488002,-487999,-487997,-487994,-487992,-487989,-487987,-487984,-487982,-487979,-487977,-487974,-487972,-487969,-487967,-487964,-487962,-487959,-487957,-487954,-487952,-487949,-487947,-487944,-487942,-487939,-487937,-487934,-487932,-487929,-487927,-487924,-487922,-487919,-487917,-487915,-487912,-487910,-487907,-487905,-487902,-487900,-487897,-487895,-487892,-487890,-487887,-487885,-487882,-487880,-487877,-487875,-487872,-487870,-487867,-487865,-487862,-487860,-487857,-487855,-487852,-487850,-487847,-487845,-487842,-487840,-487837,-487835,-487832,-487830,-487827,-487825,-487822,-487820,-487817,-487815,-487812,-487810,-487807,-487805,-487802,-487800,-487797,-487795,-487792,-487790,-487787,-487785,-487782,-487780,-487777,-487775,-487772,-487770,-487767,-487765,-487762,-487760,-487757,-487755,-487752,-487750,-487747,-487745,-487742,-487740,-487737,-487735,-487732,-487730,-487727,-487725,-487722,-487720,-487717,-487715,-487712,-487710,-487707,-487705,-487702,-487700,-487697,-487695,-487692,-487690,-487687,-487685,-487682,-487680,-487677,-487675,-487672,-487670,-487667,-487665,-487662,-487660,-487657,-487655,-487652,-487650,-487647,-487645,-487642,-487640,-487637,-487635,-487632,-487630,-487627,-487625,-487622,-487620,-487617,-487615,-487612,-487610,-487607,-487605,-487602,-487600,-487597,-487595,-487592,-487590,-487587,-487585,-487582,-487580,-487577,-487575,-487572,-487570,-487567,-487565,-487562,-487560,-487557,-487555,-487552,-487550,-487547,-487545,-487542,-487540,-487537,-487535,-487532,-487530,-487527,-487525,-487522,-487520,-487517,-487515,-487512,-487510,-487507,-487504,-487502,-487499,-487497,-487494,-487492,-487489,-487487,-487484,-487482,-487479,-487477,-487474,-487472,-487469,-487467,-487464,-487462,-487459,-487457,-487454,-487452,-487449,-487447,-487444,-487442,-487439,-487437,-487434,-487432,-487429,-487427,-487424,-487422,-487419,-487417,-487414,-487412,-487409,-487406,-487404,-487401,-487399,-487396,-487394,-487391,-487389,-487386,-487384,-487381,-487379,-487376,-487374,-487371,-487369,-487366,-487364,-487361,-487359,-487356,-487354,-487351,-487349,-487346,-487344,-487341,-487339,-487336,-487333,-487331,-487328,-487326,-487323,-487321,-487318,-487316,-487313,-487311,-487308,-487306,-487303,-487301,-487298,-487296,-487293,-487291,-487288,-487286,-487283,-487281,-487278,-487275,-487273,-487270,-487268,-487265,-487263,-487260,-487258,-487255,-487253,-487250,-487248,-487245,-487243,-487240,-487238,-487235,-487233,-487230,-487228,-487225,-487222,-487220,-487217,-487215,-487212,-487210,-487207,-487205,-487202,-487200,-487197,-487195,-487192,-487190,-487187,-487185,-487182,-487180,-487177,-487174,-487172,-487169,-487167,-487164,-487162,-487159,-487157,-487154,-487152,-487149,-487147,-487144,-487142,-487139,-487137,-487134,-487131,-487129,-487126,-487124,-487121,-487119,-487116,-487114,-487111,-487109,-487106,-487104,-487101,-487099,-487096,-487094,-487091,-487088,-487086,-487083,-487081,-487078,-487076,-487073,-487071,-487068,-487066,-487063,-487061,-487058,-487056,-487053,-487050,-487048,-487045,-487043,-487040,-487038,-487035,-487033,-487030,-487028,-487025,-487023,-487020,-487017,-487015,-487012,-487010,-487007,-487005,-487002,-487000,-486997,-486995,-486992,-486990,-486987,-486985,-486982,-486979,-486977,-486974,-486972,-486969,-486967,-486964,-486962,-486959,-486957,-486954,-486952,-486949,-486946,-486944,-486941,-486939,-486936,-486934,-486931,-486929,-486926,-486924,-486921,-486918,-486916,-486913,-486911,-486908,-486906,-486903,-486901,-486898,-486896,-486893,-486891,-486888,-486885,-486883,-486880,-486878,-486875,-486873,-486870,-486868,-486865,-486863,-486860,-486857,-486855,-486852,-486850,-486847,-486845,-486842,-486840,-486837,-486835,-486832,-486829,-486827,-486824,-486822,-486819,-486817,-486814,-486812,-486809,-486807,-486804,-486801,-486799,-486796,-486794,-486791,-486789,-486786,-486784,-486781,-486779,-486776,-486773,-486771,-486768,-486766,-486763,-486761,-486758,-486756,-486753,-486750,-486748,-486745,-486743,-486740,-486738,-486735,-486733,-486730,-486728,-486725,-486722,-486720,-486717,-486715,-486712,-486710,-486707,-486705,-486702,-486699,-486697,-486694,-486692,-486689,-486687,-486684,-486682,-486679,-486676,-486674,-486671,-486669,-486666,-486664,-486661,-486659,-486656,-486654,-486651,-486648,-486646,-486643,-486641,-486638,-486636,-486633,-486631,-486628,-486625,-486623,-486620,-486618,-486615,-486613,-486610,-486607,-486605,-486602,-486600,-486597,-486595,-486592,-486590,-486587,-486584,-486582,-486579,-486577,-486574,-486572,-486569,-486567,-486564,-486561,-486559,-486556,-486554,-486551,-486549,-486546,-486544,-486541,-486538,-486536,-486533,-486531,-486528,-486526,-486523,-486520,-486518,-486515,-486513,-486510,-486508,-486505,-486503,-486500,-486497,-486495,-486492,-486490,-486487,-486485,-486482,-486479,-486477,-486474,-486472,-486469,-486467,-486464,-486462,-486459,-486456,-486454,-486451,-486449,-486446,-486444,-486441,-486438,-486436,-486433,-486431,-486428,-486426,-486423,-486420,-486418,-486415,-486413,-486410,-486408,-486405,-486403,-486400,-486397,-486395,-486392,-486390,-486387,-486385,-486382,-486379,-486377,-486374,-486372,-486369,-486367,-486364,-486361,-486359,-486356,-486354,-486351,-486349,-486346,-486343,-486341,-486338,-486336,-486333,-486331,-486328,-486325,-486323,-486320,-486318,-486315,-486313,-486310,-486307,-486305,-486302,-486300,-486297,-486295,-486292,-486289,-486287,-486284,-486282,-486279,-486277,-486274,-486271,-486269,-486266,-486264,-486261,-486259,-486256,-486253,-486251,-486248,-486246,-486243,-486241,-486238,-486235,-486233,-486230,-486228,-486225,-486222,-486220,-486217,-486215,-486212,-486210,-486207,-486204,-486202,-486199,-486197,-486194,-486192,-486189,-486186,-486184,-486181,-486179,-486176,-486174,-486171,-486168,-486166,-486163,-486161,-486158,-486155,-486153,-486150,-486148,-486145,-486143,-486140,-486137,-486135,-486132,-486130,-486127,-486124,-486122,-486119,-486117,-486114,-486112,-486109,-486106,-486104,-486101,-486099,-486096,-486093,-486091,-486088,-486086,-486083,-486081,-486078,-486075,-486073,-486070,-486068,-486065,-486062,-486060,-486057,-486055,-486052,-486050,-486047,-486044,-486042,-486039,-486037,-486034,-486031,-486029,-486026,-486024,-486021,-486019,-486016,-486013,-486011,-486008,-486006,-486003,-486000,-485998,-485995,-485993,-485990,-485987,-485985,-485982,-485980,-485977,-485975,-485972,-485969,-485967,-485964,-485962,-485959,-485956,-485954,-485951,-485949,-485946,-485943,-485941,-485938,-485936,-485933,-485931,-485928,-485925,-485923,-485920,-485918,-485915,-485912,-485910,-485907,-485905,-485902,-485899,-485897,-485894,-485892,-485889,-485886,-485884,-485881,-485879,-485876,-485873,-485871,-485868,-485866,-485863,-485861,-485858,-485855,-485853,-485850,-485848,-485845,-485842,-485840,-485837,-485835,-485832,-485829,-485827,-485824,-485822,-485819,-485816,-485814,-485811,-485809,-485806,-485803,-485801,-485798,-485796,-485793,-485790,-485788,-485785,-485783,-485780,-485777,-485775,-485772,-485770,-485767,-485764,-485762,-485759,-485757,-485754,-485751,-485749,-485746,-485744,-485741,-485738,-485736,-485733,-485731,-485728,-485725,-485723,-485720,-485718,-485715,-485712,-485710,-485707,-485705,-485702,-485699,-485697,-485694,-485692,-485689,-485686,-485684,-485681,-485679,-485676,-485673,-485671,-485668,-485666,-485663,-485660,-485658,-485655,-485653,-485650,-485647,-485645,-485642,-485639,-485637,-485634,-485632,-485629,-485626,-485624,-485621,-485619,-485616,-485613,-485611,-485608,-485606,-485603,-485600,-485598,-485595,-485593,-485590,-485587,-485585,-485582,-485580,-485577,-485574,-485572,-485569,-485566,-485564,-485561,-485559,-485556,-485553,-485551,-485548,-485546,-485543,-485540,-485538,-485535,-485533,-485530,-485527,-485525,-485522,-485519,-485517,-485514,-485512,-485509,-485506,-485504,-485501,-485499,-485496,-485493,-485491,-485488,-485486,-485483,-485480,-485478,-485475,-485472,-485470,-485467,-485465,-485462,-485459,-485457,-485454,-485452,-485449,-485446,-485444,-485441,-485438,-485436,-485433,-485431,-485428,-485425,-485423,-485420,-485418,-485415,-485412,-485410,-485407,-485404,-485402,-485399,-485397,-485394,-485391,-485389,-485386,-485383,-485381,-485378,-485376,-485373,-485370,-485368,-485365,-485363,-485360,-485357,-485355,-485352,-485349,-485347,-485344,-485342,-485339,-485336,-485334,-485331,-485328,-485326,-485323,-485321,-485318,-485315,-485313,-485310,-485307,-485305,-485302,-485300,-485297,-485294,-485292,-485289,-485287,-485284,-485281,-485279,-485276,-485273,-485271,-485268,-485266,-485263,-485260,-485258,-485255,-485252,-485250,-485247,-485245,-485242,-485239,-485237,-485234,-485231,-485229,-485226,-485224,-485221,-485218,-485216,-485213,-485210,-485208,-485205,-485203,-485200,-485197,-485195,-485192,-485189,-485187,-485184,-485181,-485179,-485176,-485174,-485171,-485168,-485166,-485163,-485160,-485158,-485155,-485153,-485150,-485147,-485145,-485142,-485139,-485137,-485134,-485132,-485129,-485126,-485124,-485121,-485118,-485116,-485113,-485110,-485108,-485105,-485103,-485100,-485097,-485095,-485092,-485089,-485087,-485084,-485082,-485079,-485076,-485074,-485071,-485068,-485066,-485063,-485060,-485058,-485055,-485053,-485050,-485047,-485045,-485042,-485039,-485037,-485034,-485031,-485029,-485026,-485024,-485021,-485018,-485016,-485013,-485010,-485008,-485005,-485002,-485000,-484997,-484995,-484992,-484989,-484987,-484984,-484981,-484979,-484976,-484973,-484971,-484968,-484966,-484963,-484960,-484958,-484955,-484952,-484950,-484947,-484944,-484942,-484939,-484936,-484934,-484931,-484929,-484926,-484923,-484921,-484918,-484915,-484913,-484910,-484907,-484905,-484902,-484899,-484897,-484894,-484892,-484889,-484886,-484884,-484881,-484878,-484876,-484873,-484870,-484868,-484865,-484862,-484860,-484857,-484855,-484852,-484849,-484847,-484844,-484841,-484839,-484836,-484833,-484831,-484828,-484825,-484823,-484820,-484818,-484815,-484812,-484810,-484807,-484804,-484802,-484799,-484796,-484794,-484791,-484788,-484786,-484783,-484780,-484778,-484775,-484772,-484770,-484767,-484765,-484762,-484759,-484757,-484754,-484751,-484749,-484746,-484743,-484741,-484738,-484735,-484733,-484730,-484727,-484725,-484722,-484719,-484717,-484714,-484712,-484709,-484706,-484704,-484701,-484698,-484696,-484693,-484690,-484688,-484685,-484682,-484680,-484677,-484674,-484672,-484669,-484666,-484664,-484661,-484658,-484656,-484653,-484651,-484648,-484645,-484643,-484640,-484637,-484635,-484632,-484629,-484627,-484624,-484621,-484619,-484616,-484613,-484611,-484608,-484605,-484603,-484600,-484597,-484595,-484592,-484589,-484587,-484584,-484581,-484579,-484576,-484573,-484571,-484568,-484566,-484563,-484560,-484558,-484555,-484552,-484550,-484547,-484544,-484542,-484539,-484536,-484534,-484531,-484528,-484526,-484523,-484520,-484518,-484515,-484512,-484510,-484507,-484504,-484502,-484499,-484496,-484494,-484491,-484488,-484486,-484483,-484480,-484478,-484475,-484472,-484470,-484467,-484464,-484462,-484459,-484456,-484454,-484451,-484448,-484446,-484443,-484440,-484438,-484435,-484432,-484430,-484427,-484424,-484422,-484419,-484416,-484414,-484411,-484408,-484406,-484403,-484400,-484398,-484395,-484392,-484390,-484387,-484384,-484382,-484379,-484376,-484374,-484371,-484368,-484366,-484363,-484360,-484358,-484355,-484352,-484350,-484347,-484344,-484342,-484339,-484336,-484334,-484331,-484328,-484326,-484323,-484320,-484318,-484315,-484312,-484310,-484307,-484304,-484302,-484299,-484296,-484294,-484291,-484288,-484286,-484283,-484280,-484278,-484275,-484272,-484270,-484267,-484264,-484262,-484259,-484256,-484254,-484251,-484248,-484246,-484243,-484240,-484237,-484235,-484232,-484229,-484227,-484224,-484221,-484219,-484216,-484213,-484211,-484208,-484205,-484203,-484200,-484197,-484195,-484192,-484189,-484187,-484184,-484181,-484179,-484176,-484173,-484171,-484168,-484165,-484163,-484160,-484157,-484155,-484152,-484149,-484146,-484144,-484141,-484138,-484136,-484133,-484130,-484128,-484125,-484122,-484120,-484117,-484114,-484112,-484109,-484106,-484104,-484101,-484098,-484096,-484093,-484090,-484088,-484085,-484082,-484079,-484077,-484074,-484071,-484069,-484066,-484063,-484061,-484058,-484055,-484053,-484050,-484047,-484045,-484042,-484039,-484037,-484034,-484031,-484028,-484026,-484023,-484020,-484018,-484015,-484012,-484010,-484007,-484004,-484002,-483999,-483996,-483994,-483991,-483988,-483986,-483983,-483980,-483977,-483975,-483972,-483969,-483967,-483964,-483961,-483959,-483956,-483953,-483951,-483948,-483945,-483942,-483940,-483937,-483934,-483932,-483929,-483926,-483924,-483921,-483918,-483916,-483913,-483910,-483908,-483905,-483902,-483899,-483897,-483894,-483891,-483889,-483886,-483883,-483881,-483878,-483875,-483873,-483870,-483867,-483864,-483862,-483859,-483856,-483854,-483851,-483848,-483846,-483843,-483840,-483838,-483835,-483832,-483829,-483827,-483824,-483821,-483819,-483816,-483813,-483811,-483808,-483805,-483802,-483800,-483797,-483794,-483792,-483789,-483786,-483784,-483781,-483778,-483776,-483773,-483770,-483767,-483765,-483762,-483759,-483757,-483754,-483751,-483749,-483746,-483743,-483740,-483738,-483735,-483732,-483730,-483727,-483724,-483722,-483719,-483716,-483713,-483711,-483708,-483705,-483703,-483700,-483697,-483695,-483692,-483689,-483686,-483684,-483681,-483678,-483676,-483673,-483670,-483668,-483665,-483662,-483659,-483657,-483654,-483651,-483649,-483646,-483643,-483641,-483638,-483635,-483632,-483630,-483627,-483624,-483622,-483619,-483616,-483613,-483611,-483608,-483605,-483603,-483600,-483597,-483595,-483592,-483589,-483586,-483584,-483581,-483578,-483576,-483573,-483570,-483567,-483565,-483562,-483559,-483557,-483554,-483551,-483549,-483546,-483543,-483540,-483538,-483535,-483532,-483530,-483527,-483524,-483521,-483519,-483516,-483513,-483511,-483508,-483505,-483502,-483500,-483497,-483494,-483492,-483489,-483486,-483483,-483481,-483478,-483475,-483473,-483470,-483467,-483465,-483462,-483459,-483456,-483454,-483451,-483448,-483446,-483443,-483440,-483437,-483435,-483432,-483429,-483427,-483424,-483421,-483418,-483416,-483413,-483410,-483408,-483405,-483402,-483399,-483397,-483394,-483391,-483389,-483386,-483383,-483380,-483378,-483375,-483372,-483370,-483367,-483364,-483361,-483359,-483356,-483353,-483351,-483348,-483345,-483342,-483340,-483337,-483334,-483331,-483329,-483326,-483323,-483321,-483318,-483315,-483312,-483310,-483307,-483304,-483302,-483299,-483296,-483293,-483291,-483288,-483285,-483283,-483280,-483277,-483274,-483272,-483269,-483266,-483263,-483261,-483258,-483255,-483253,-483250,-483247,-483244,-483242,-483239,-483236,-483234,-483231,-483228,-483225,-483223,-483220,-483217,-483214,-483212,-483209,-483206,-483204,-483201,-483198,-483195,-483193,-483190,-483187,-483185,-483182,-483179,-483176,-483174,-483171,-483168,-483165,-483163,-483160,-483157,-483155,-483152,-483149,-483146,-483144,-483141,-483138,-483135,-483133,-483130,-483127,-483125,-483122,-483119,-483116,-483114,-483111,-483108,-483105,-483103,-483100,-483097,-483095,-483092,-483089,-483086,-483084,-483081,-483078,-483075,-483073,-483070,-483067,-483064,-483062,-483059,-483056,-483054,-483051,-483048,-483045,-483043,-483040,-483037,-483034,-483032,-483029,-483026,-483023,-483021,-483018,-483015,-483013,-483010,-483007,-483004,-483002,-482999,-482996,-482993,-482991,-482988,-482985,-482982,-482980,-482977,-482974,-482972,-482969,-482966,-482963,-482961,-482958,-482955,-482952,-482950,-482947,-482944,-482941,-482939,-482936,-482933,-482930,-482928,-482925,-482922,-482920,-482917,-482914,-482911,-482909,-482906,-482903,-482900,-482898,-482895,-482892,-482889,-482887,-482884,-482881,-482878,-482876,-482873,-482870,-482868,-482865,-482862,-482859,-482857,-482854,-482851,-482848,-482846,-482843,-482840,-482837,-482835,-482832,-482829,-482826,-482824,-482821,-482818,-482815,-482813,-482810,-482807,-482804,-482802,-482799,-482796,-482793,-482791,-482788,-482785,-482782,-482780,-482777,-482774,-482772,-482769,-482766,-482763,-482761,-482758,-482755,-482752,-482750,-482747,-482744,-482741,-482739,-482736,-482733,-482730,-482728,-482725,-482722,-482719,-482717,-482714,-482711,-482708,-482706,-482703,-482700,-482697,-482695,-482692,-482689,-482686,-482684,-482681,-482678,-482675,-482673,-482670,-482667,-482664,-482662,-482659,-482656,-482653,-482651,-482648,-482645,-482642,-482640,-482637,-482634,-482631,-482629,-482626,-482623,-482620,-482618,-482615,-482612,-482609,-482607,-482604,-482601,-482598,-482596,-482593,-482590,-482587,-482585,-482582,-482579,-482576,-482574,-482571,-482568,-482565,-482563,-482560,-482557,-482554,-482552,-482549,-482546,-482543,-482541,-482538,-482535,-482532,-482529,-482527,-482524,-482521,-482518,-482516,-482513,-482510,-482507,-482505,-482502,-482499,-482496,-482494,-482491,-482488,-482485,-482483,-482480,-482477,-482474,-482472,-482469,-482466,-482463,-482461,-482458,-482455,-482452,-482450,-482447,-482444,-482441,-482438,-482436,-482433,-482430,-482427,-482425,-482422,-482419,-482416,-482414,-482411,-482408,-482405,-482403,-482400,-482397,-482394,-482392,-482389,-482386,-482383,-482380,-482378,-482375,-482372,-482369,-482367,-482364,-482361,-482358,-482356,-482353,-482350,-482347,-482345,-482342,-482339,-482336,-482333,-482331,-482328,-482325,-482322,-482320,-482317,-482314,-482311,-482309,-482306,-482303,-482300,-482298,-482295,-482292,-482289,-482286,-482284,-482281,-482278,-482275,-482273,-482270,-482267,-482264,-482262,-482259,-482256,-482253,-482250,-482248,-482245,-482242,-482239,-482237,-482234,-482231,-482228,-482226,-482223,-482220,-482217,-482214,-482212,-482209,-482206,-482203,-482201,-482198,-482195,-482192,-482190,-482187,-482184,-482181,-482178,-482176,-482173,-482170,-482167,-482165,-482162,-482159,-482156,-482153,-482151,-482148,-482145,-482142,-482140,-482137,-482134,-482131,-482128,-482126,-482123,-482120,-482117,-482115,-482112,-482109,-482106,-482104,-482101,-482098,-482095,-482092,-482090,-482087,-482084,-482081,-482079,-482076,-482073,-482070,-482067,-482065,-482062,-482059,-482056,-482054,-482051,-482048,-482045,-482042,-482040,-482037,-482034,-482031,-482029,-482026,-482023,-482020,-482017,-482015,-482012,-482009,-482006,-482003,-482001,-481998,-481995,-481992,-481990,-481987,-481984,-481981,-481978,-481976,-481973,-481970,-481967,-481965,-481962,-481959,-481956,-481953,-481951,-481948,-481945,-481942,-481939,-481937,-481934,-481931,-481928,-481926,-481923,-481920,-481917,-481914,-481912,-481909,-481906,-481903,-481901,-481898,-481895,-481892,-481889,-481887,-481884,-481881,-481878,-481875,-481873,-481870,-481867,-481864,-481862,-481859,-481856,-481853,-481850,-481848,-481845,-481842,-481839,-481836,-481834,-481831,-481828,-481825,-481822,-481820,-481817,-481814,-481811,-481809,-481806,-481803,-481800,-481797,-481795,-481792,-481789,-481786,-481783,-481781,-481778,-481775,-481772,-481769,-481767,-481764,-481761,-481758,-481755,-481753,-481750,-481747,-481744,-481742,-481739,-481736,-481733,-481730,-481728,-481725,-481722,-481719,-481716,-481714,-481711,-481708,-481705,-481702,-481700,-481697,-481694,-481691,-481688,-481686,-481683,-481680,-481677,-481674,-481672,-481669,-481666,-481663,-481660,-481658,-481655,-481652,-481649,-481647,-481644,-481641,-481638,-481635,-481633,-481630,-481627,-481624,-481621,-481619,-481616,-481613,-481610,-481607,-481605,-481602,-481599,-481596,-481593,-481591,-481588,-481585,-481582,-481579,-481577,-481574,-481571,-481568,-481565,-481563,-481560,-481557,-481554,-481551,-481549,-481546,-481543,-481540,-481537,-481535,-481532,-481529,-481526,-481523,-481521,-481518,-481515,-481512,-481509,-481506,-481504,-481501,-481498,-481495,-481492,-481490,-481487,-481484,-481481,-481478,-481476,-481473,-481470,-481467,-481464,-481462,-481459,-481456,-481453,-481450,-481448,-481445,-481442,-481439,-481436,-481434,-481431,-481428,-481425,-481422,-481420,-481417,-481414,-481411,-481408,-481405,-481403,-481400,-481397,-481394,-481391,-481389,-481386,-481383,-481380,-481377,-481375,-481372,-481369,-481366,-481363,-481361,-481358,-481355,-481352,-481349,-481346,-481344,-481341,-481338,-481335,-481332,-481330,-481327,-481324,-481321,-481318,-481316,-481313,-481310,-481307,-481304,-481301,-481299,-481296,-481293,-481290,-481287,-481285,-481282,-481279,-481276,-481273,-481271,-481268,-481265,-481262,-481259,-481256,-481254,-481251,-481248,-481245,-481242,-481240,-481237,-481234,-481231,-481228,-481225,-481223,-481220,-481217,-481214,-481211,-481209,-481206,-481203,-481200,-481197,-481194,-481192,-481189,-481186,-481183,-481180,-481178,-481175,-481172,-481169,-481166,-481163,-481161,-481158,-481155,-481152,-481149,-481147,-481144,-481141,-481138,-481135,-481132,-481130,-481127,-481124,-481121,-481118,-481116,-481113,-481110,-481107,-481104,-481101,-481099,-481096,-481093,-481090,-481087,-481084,-481082,-481079,-481076,-481073,-481070,-481068,-481065,-481062,-481059,-481056,-481053,-481051,-481048,-481045,-481042,-481039,-481036,-481034,-481031,-481028,-481025,-481022,-481020,-481017,-481014,-481011,-481008,-481005,-481003,-481000,-480997,-480994,-480991,-480988,-480986,-480983,-480980,-480977,-480974,-480971,-480969,-480966,-480963,-480960,-480957,-480955,-480952,-480949,-480946,-480943,-480940,-480938,-480935,-480932,-480929,-480926,-480923,-480921,-480918,-480915,-480912,-480909,-480906,-480904,-480901,-480898,-480895,-480892,-480889,-480887,-480884,-480881,-480878,-480875,-480872,-480870,-480867,-480864,-480861,-480858,-480855,-480853,-480850,-480847,-480844,-480841,-480838,-480836,-480833,-480830,-480827,-480824,-480821,-480819,-480816,-480813,-480810,-480807,-480804,-480802,-480799,-480796,-480793,-480790,-480787,-480785,-480782,-480779,-480776,-480773,-480770,-480768,-480765,-480762,-480759,-480756,-480753,-480750,-480748,-480745,-480742,-480739,-480736,-480733,-480731,-480728,-480725,-480722,-480719,-480716,-480714,-480711,-480708,-480705,-480702,-480699,-480697,-480694,-480691,-480688,-480685,-480682,-480679,-480677,-480674,-480671,-480668,-480665,-480662,-480660,-480657,-480654,-480651,-480648,-480645,-480643,-480640,-480637,-480634,-480631,-480628,-480625,-480623,-480620,-480617,-480614,-480611,-480608,-480606,-480603,-480600,-480597,-480594,-480591,-480589,-480586,-480583,-480580,-480577,-480574,-480571,-480569,-480566,-480563,-480560,-480557,-480554,-480552,-480549,-480546,-480543,-480540,-480537,-480534,-480532,-480529,-480526,-480523,-480520,-480517,-480514,-480512,-480509,-480506,-480503,-480500,-480497,-480495,-480492,-480489,-480486,-480483,-480480,-480477,-480475,-480472,-480469,-480466,-480463,-480460,-480457,-480455,-480452,-480449,-480446,-480443,-480440,-480438,-480435,-480432,-480429,-480426,-480423,-480420,-480418,-480415,-480412,-480409,-480406,-480403,-480400,-480398,-480395,-480392,-480389,-480386,-480383,-480380,-480378,-480375,-480372,-480369,-480366,-480363,-480360,-480358,-480355,-480352,-480349,-480346,-480343,-480340,-480338,-480335,-480332,-480329,-480326,-480323,-480320,-480318,-480315,-480312,-480309,-480306,-480303,-480300,-480298,-480295,-480292,-480289,-480286,-480283,-480280,-480278,-480275,-480272,-480269,-480266,-480263,-480260,-480258,-480255,-480252,-480249,-480246,-480243,-480240,-480238,-480235,-480232,-480229,-480226,-480223,-480220,-480218,-480215,-480212,-480209,-480206,-480203,-480200,-480197,-480195,-480192,-480189,-480186,-480183,-480180,-480177,-480175,-480172,-480169,-480166,-480163,-480160,-480157,-480155,-480152,-480149,-480146,-480143,-480140,-480137,-480134,-480132,-480129,-480126,-480123,-480120,-480117,-480114,-480112,-480109,-480106,-480103,-480100,-480097,-480094,-480091,-480089,-480086,-480083,-480080,-480077,-480074,-480071,-480069,-480066,-480063,-480060,-480057,-480054,-480051,-480048,-480046,-480043,-480040,-480037,-480034,-480031,-480028,-480025,-480023,-480020,-480017,-480014,-480011,-480008,-480005,-480002,-480000,-479997,-479994,-479991,-479988,-479985,-479982,-479980,-479977,-479974,-479971,-479968,-479965,-479962,-479959,-479957,-479954,-479951,-479948,-479945,-479942,-479939,-479936,-479934,-479931,-479928,-479925,-479922,-479919,-479916,-479913,-479911,-479908,-479905,-479902,-479899,-479896,-479893,-479890,-479888,-479885,-479882,-479879,-479876,-479873,-479870,-479867,-479864,-479862,-479859,-479856,-479853,-479850,-479847,-479844,-479841,-479839,-479836,-479833,-479830,-479827,-479824,-479821,-479818,-479816,-479813,-479810,-479807,-479804,-479801,-479798,-479795,-479792,-479790,-479787,-479784,-479781,-479778,-479775,-479772,-479769,-479767,-479764,-479761,-479758,-479755,-479752,-479749,-479746,-479743,-479741,-479738,-479735,-479732,-479729,-479726,-479723,-479720,-479718,-479715,-479712,-479709,-479706,-479703,-479700,-479697,-479694,-479692,-479689,-479686,-479683,-479680,-479677,-479674,-479671,-479668,-479666,-479663,-479660,-479657,-479654,-479651,-479648,-479645,-479643,-479640,-479637,-479634,-479631,-479628,-479625,-479622,-479619,-479617,-479614,-479611,-479608,-479605,-479602,-479599,-479596,-479593,-479590,-479588,-479585,-479582,-479579,-479576,-479573,-479570,-479567,-479564,-479562,-479559,-479556,-479553,-479550,-479547,-479544,-479541,-479538,-479536,-479533,-479530,-479527,-479524,-479521,-479518,-479515,-479512,-479510,-479507,-479504,-479501,-479498,-479495,-479492,-479489,-479486,-479483,-479481,-479478,-479475,-479472,-479469,-479466,-479463,-479460,-479457,-479455,-479452,-479449,-479446,-479443,-479440,-479437,-479434,-479431,-479428,-479426,-479423,-479420,-479417,-479414,-479411,-479408,-479405,-479402,-479399,-479397,-479394,-479391,-479388,-479385,-479382,-479379,-479376,-479373,-479370,-479368,-479365,-479362,-479359,-479356,-479353,-479350,-479347,-479344,-479341,-479339,-479336,-479333,-479330,-479327,-479324,-479321,-479318,-479315,-479312,-479310,-479307,-479304,-479301,-479298,-479295,-479292,-479289,-479286,-479283,-479281,-479278,-479275,-479272,-479269,-479266,-479263,-479260,-479257,-479254,-479251,-479249,-479246,-479243,-479240,-479237,-479234,-479231,-479228,-479225,-479222,-479220,-479217,-479214,-479211,-479208,-479205,-479202,-479199,-479196,-479193,-479190,-479188,-479185,-479182,-479179,-479176,-479173,-479170,-479167,-479164,-479161,-479158,-479156,-479153,-479150,-479147,-479144,-479141,-479138,-479135,-479132,-479129,-479126,-479124,-479121,-479118,-479115,-479112,-479109,-479106,-479103,-479100,-479097,-479094,-479091,-479089,-479086,-479083,-479080,-479077,-479074,-479071,-479068,-479065,-479062,-479059,-479057,-479054,-479051,-479048,-479045,-479042,-479039,-479036,-479033,-479030,-479027,-479024,-479022,-479019,-479016,-479013,-479010,-479007,-479004,-479001,-478998,-478995,-478992,-478989,-478987,-478984,-478981,-478978,-478975,-478972,-478969,-478966,-478963,-478960,-478957,-478954,-478952,-478949,-478946,-478943,-478940,-478937,-478934,-478931,-478928,-478925,-478922,-478919,-478917,-478914,-478911,-478908,-478905,-478902,-478899,-478896,-478893,-478890,-478887,-478884,-478881,-478879,-478876,-478873,-478870,-478867,-478864,-478861,-478858,-478855,-478852,-478849,-478846,-478843,-478841,-478838,-478835,-478832,-478829,-478826,-478823,-478820,-478817,-478814,-478811,-478808,-478805,-478803,-478800,-478797,-478794,-478791,-478788,-478785,-478782,-478779,-478776,-478773,-478770,-478767,-478765,-478762,-478759,-478756,-478753,-478750,-478747,-478744,-478741,-478738,-478735,-478732,-478729,-478726,-478724,-478721,-478718,-478715,-478712,-478709,-478706,-478703,-478700,-478697,-478694,-478691,-478688,-478685,-478683,-478680,-478677,-478674,-478671,-478668,-478665,-478662,-478659,-478656,-478653,-478650,-478647,-478644,-478641,-478639,-478636,-478633,-478630,-478627,-478624,-478621,-478618,-478615,-478612,-478609,-478606,-478603,-478600,-478597,-478595,-478592,-478589,-478586,-478583,-478580,-478577,-478574,-478571,-478568,-478565,-478562,-478559,-478556,-478553,-478551,-478548,-478545,-478542,-478539,-478536,-478533,-478530,-478527,-478524,-478521,-478518,-478515,-478512,-478509,-478506,-478504,-478501,-478498,-478495,-478492,-478489,-478486,-478483,-478480,-478477,-478474,-478471,-478468,-478465,-478462,-478459,-478457,-478454,-478451,-478448,-478445,-478442,-478439,-478436,-478433,-478430,-478427,-478424,-478421,-478418,-478415,-478412,-478409,-478407,-478404,-478401,-478398,-478395,-478392,-478389,-478386,-478383,-478380,-478377,-478374,-478371,-478368,-478365,-478362,-478359,-478356,-478354,-478351,-478348,-478345,-478342,-478339,-478336,-478333,-478330,-478327,-478324,-478321,-478318,-478315,-478312,-478309,-478306,-478303,-478300,-478298,-478295,-478292,-478289,-478286,-478283,-478280,-478277,-478274,-478271,-478268,-478265,-478262,-478259,-478256,-478253,-478250,-478247,-478244,-478242,-478239,-478236,-478233,-478230,-478227,-478224,-478221,-478218,-478215,-478212,-478209,-478206,-478203,-478200,-478197,-478194,-478191,-478188,-478185,-478183,-478180,-478177,-478174,-478171,-478168,-478165,-478162,-478159,-478156,-478153,-478150,-478147,-478144,-478141,-478138,-478135,-478132,-478129,-478126,-478123,-478121,-478118,-478115,-478112,-478109,-478106,-478103,-478100,-478097,-478094,-478091,-478088,-478085,-478082,-478079,-478076,-478073,-478070,-478067,-478064,-478061,-478058,-478055,-478053,-478050,-478047,-478044,-478041,-478038,-478035,-478032,-478029,-478026,-478023,-478020,-478017,-478014,-478011,-478008,-478005,-478002,-477999,-477996,-477993,-477990,-477987,-477984,-477981,-477979,-477976,-477973,-477970,-477967,-477964,-477961,-477958,-477955,-477952,-477949,-477946,-477943,-477940,-477937,-477934,-477931,-477928,-477925,-477922,-477919,-477916,-477913,-477910,-477907,-477904,-477902,-477899,-477896,-477893,-477890,-477887,-477884,-477881,-477878,-477875,-477872,-477869,-477866,-477863,-477860,-477857,-477854,-477851,-477848,-477845,-477842,-477839,-477836,-477833,-477830,-477827,-477824,-477821,-477818,-477815,-477813,-477810,-477807,-477804,-477801,-477798,-477795,-477792,-477789,-477786,-477783,-477780,-477777,-477774,-477771,-477768,-477765,-477762,-477759,-477756,-477753,-477750,-477747,-477744,-477741,-477738,-477735,-477732,-477729,-477726,-477723,-477720,-477717,-477715,-477712,-477709,-477706,-477703,-477700,-477697,-477694,-477691,-477688,-477685,-477682,-477679,-477676,-477673,-477670,-477667,-477664,-477661,-477658,-477655,-477652,-477649,-477646,-477643,-477640,-477637,-477634,-477631,-477628,-477625,-477622,-477619,-477616,-477613,-477610,-477607,-477604,-477601,-477598,-477596,-477593,-477590,-477587,-477584,-477581,-477578,-477575,-477572,-477569,-477566,-477563,-477560,-477557,-477554,-477551,-477548,-477545,-477542,-477539,-477536,-477533,-477530,-477527,-477524,-477521,-477518,-477515,-477512,-477509,-477506,-477503,-477500,-477497,-477494,-477491,-477488,-477485,-477482,-477479,-477476,-477473,-477470,-477467,-477464,-477461,-477458,-477455,-477452,-477449,-477446,-477444,-477441,-477438,-477435,-477432,-477429,-477426,-477423,-477420,-477417,-477414,-477411,-477408,-477405,-477402,-477399,-477396,-477393,-477390,-477387,-477384,-477381,-477378,-477375,-477372,-477369,-477366,-477363,-477360,-477357,-477354,-477351,-477348,-477345,-477342,-477339,-477336,-477333,-477330,-477327,-477324,-477321,-477318,-477315,-477312,-477309,-477306,-477303,-477300,-477297,-477294,-477291,-477288,-477285,-477282,-477279,-477276,-477273,-477270,-477267,-477264,-477261,-477258,-477255,-477252,-477249,-477246,-477243,-477240,-477237,-477234,-477231,-477228,-477225,-477222,-477219,-477216,-477213,-477210,-477207,-477204,-477201,-477198,-477195,-477192,-477189,-477186,-477183,-477180,-477177,-477174,-477171,-477168,-477165,-477162,-477159,-477156,-477153,-477150,-477147,-477144,-477141,-477138,-477135,-477132,-477129,-477126,-477124,-477121,-477118,-477115,-477112,-477109,-477106,-477103,-477100,-477097,-477094,-477091,-477088,-477085,-477082,-477079,-477076,-477073,-477070,-477067,-477064,-477061,-477058,-477055,-477052,-477049,-477046,-477043,-477040,-477037,-477034,-477031,-477028,-477025,-477022,-477019,-477016,-477013,-477010,-477007,-477003,-477000,-476997,-476994,-476991,-476988,-476985,-476982,-476979,-476976,-476973,-476970,-476967,-476964,-476961,-476958,-476955,-476952,-476949,-476946,-476943,-476940,-476937,-476934,-476931,-476928,-476925,-476922,-476919,-476916,-476913,-476910,-476907,-476904,-476901,-476898,-476895,-476892,-476889,-476886,-476883,-476880,-476877,-476874,-476871,-476868,-476865,-476862,-476859,-476856,-476853,-476850,-476847,-476844,-476841,-476838,-476835,-476832,-476829,-476826,-476823,-476820,-476817,-476814,-476811,-476808,-476805,-476802,-476799,-476796,-476793,-476790,-476787,-476784,-476781,-476778,-476775,-476772,-476769,-476766,-476763,-476760,-476757,-476754,-476751,-476748,-476745,-476742,-476739,-476736,-476733,-476730,-476727,-476724,-476721,-476718,-476715,-476712,-476709,-476706,-476703,-476700,-476697,-476694,-476691,-476688,-476685,-476681,-476678,-476675,-476672,-476669,-476666,-476663,-476660,-476657,-476654,-476651,-476648,-476645,-476642,-476639,-476636,-476633,-476630,-476627,-476624,-476621,-476618,-476615,-476612,-476609,-476606,-476603,-476600,-476597,-476594,-476591,-476588,-476585,-476582,-476579,-476576,-476573,-476570,-476567,-476564,-476561,-476558,-476555,-476552,-476549,-476546,-476543,-476540,-476537,-476534,-476531,-476527,-476524,-476521,-476518,-476515,-476512,-476509,-476506,-476503,-476500,-476497,-476494,-476491,-476488,-476485,-476482,-476479,-476476,-476473,-476470,-476467,-476464,-476461,-476458,-476455,-476452,-476449,-476446,-476443,-476440,-476437,-476434,-476431,-476428,-476425,-476422,-476419,-476416,-476413,-476410,-476406,-476403,-476400,-476397,-476394,-476391,-476388,-476385,-476382,-476379,-476376,-476373,-476370,-476367,-476364,-476361,-476358,-476355,-476352,-476349,-476346,-476343,-476340,-476337,-476334,-476331,-476328,-476325,-476322,-476319,-476316,-476313,-476310,-476306,-476303,-476300,-476297,-476294,-476291,-476288,-476285,-476282,-476279,-476276,-476273,-476270,-476267,-476264,-476261,-476258,-476255,-476252,-476249,-476246,-476243,-476240,-476237,-476234,-476231,-476228,-476225,-476222,-476218,-476215,-476212,-476209,-476206,-476203,-476200,-476197,-476194,-476191,-476188,-476185,-476182,-476179,-476176,-476173,-476170,-476167,-476164,-476161,-476158,-476155,-476152,-476149,-476146,-476143,-476140,-476136,-476133,-476130,-476127,-476124,-476121,-476118,-476115,-476112,-476109,-476106,-476103,-476100,-476097,-476094,-476091,-476088,-476085,-476082,-476079,-476076,-476073,-476070,-476067,-476064,-476060,-476057,-476054,-476051,-476048,-476045,-476042,-476039,-476036,-476033,-476030,-476027,-476024,-476021,-476018,-476015,-476012,-476009,-476006,-476003,-476000,-475997,-475994,-475990,-475987,-475984,-475981,-475978,-475975,-475972,-475969,-475966,-475963,-475960,-475957,-475954,-475951,-475948,-475945,-475942,-475939,-475936,-475933,-475930,-475926,-475923,-475920,-475917,-475914,-475911,-475908,-475905,-475902,-475899,-475896,-475893,-475890,-475887,-475884,-475881,-475878,-475875,-475872,-475869,-475865,-475862,-475859,-475856,-475853,-475850,-475847,-475844,-475841,-475838,-475835,-475832,-475829,-475826,-475823,-475820,-475817,-475814,-475811,-475808,-475804,-475801,-475798,-475795,-475792,-475789,-475786,-475783,-475780,-475777,-475774,-475771,-475768,-475765,-475762,-475759,-475756,-475753,-475749,-475746,-475743,-475740,-475737,-475734,-475731,-475728,-475725,-475722,-475719,-475716,-475713,-475710,-475707,-475704,-475701,-475698,-475694,-475691,-475688,-475685,-475682,-475679,-475676,-475673,-475670,-475667,-475664,-475661,-475658,-475655,-475652,-475649,-475646,-475642,-475639,-475636,-475633,-475630,-475627,-475624,-475621,-475618,-475615,-475612,-475609,-475606,-475603,-475600,-475597,-475593,-475590,-475587,-475584,-475581,-475578,-475575,-475572,-475569,-475566,-475563,-475560,-475557,-475554,-475551,-475548,-475544,-475541,-475538,-475535,-475532,-475529,-475526,-475523,-475520,-475517,-475514,-475511,-475508,-475505,-475502,-475498,-475495,-475492,-475489,-475486,-475483,-475480,-475477,-475474,-475471,-475468,-475465,-475462,-475459,-475456,-475452,-475449,-475446,-475443,-475440,-475437,-475434,-475431,-475428,-475425,-475422,-475419,-475416,-475413,-475410,-475406,-475403,-475400,-475397,-475394,-475391,-475388,-475385,-475382,-475379,-475376,-475373,-475370,-475367,-475363,-475360,-475357,-475354,-475351,-475348,-475345,-475342,-475339,-475336,-475333,-475330,-475327,-475324,-475320,-475317,-475314,-475311,-475308,-475305,-475302,-475299,-475296,-475293,-475290,-475287,-475284,-475281,-475277,-475274,-475271,-475268,-475265,-475262,-475259,-475256,-475253,-475250,-475247,-475244,-475241,-475237,-475234,-475231,-475228,-475225,-475222,-475219,-475216,-475213,-475210,-475207,-475204,-475201,-475197,-475194,-475191,-475188,-475185,-475182,-475179,-475176,-475173,-475170,-475167,-475164,-475160,-475157,-475154,-475151,-475148,-475145,-475142,-475139,-475136,-475133,-475130,-475127,-475124,-475120,-475117,-475114,-475111,-475108,-475105,-475102,-475099,-475096,-475093,-475090,-475087,-475083,-475080,-475077,-475074,-475071,-475068,-475065,-475062,-475059,-475056,-475053,-475050,-475046,-475043,-475040,-475037,-475034,-475031,-475028,-475025,-475022,-475019,-475016,-475013,-475009,-475006,-475003,-475000,-474997,-474994,-474991,-474988,-474985,-474982,-474979,-474975,-474972,-474969,-474966,-474963,-474960,-474957,-474954,-474951,-474948,-474945,-474941,-474938,-474935,-474932,-474929,-474926,-474923,-474920,-474917,-474914,-474911,-474908,-474904,-474901,-474898,-474895,-474892,-474889,-474886,-474883,-474880,-474877,-474874,-474870,-474867,-474864,-474861,-474858,-474855,-474852,-474849,-474846,-474843,-474839,-474836,-474833,-474830,-474827,-474824,-474821,-474818,-474815,-474812,-474809,-474805,-474802,-474799,-474796,-474793,-474790,-474787,-474784,-474781,-474778,-474775,-474771,-474768,-474765,-474762,-474759,-474756,-474753,-474750,-474747,-474744,-474740,-474737,-474734,-474731,-474728,-474725,-474722,-474719,-474716,-474713,-474709,-474706,-474703,-474700,-474697,-474694,-474691,-474688,-474685,-474682,-474678,-474675,-474672,-474669,-474666,-474663,-474660,-474657,-474654,-474651,-474647,-474644,-474641,-474638,-474635,-474632,-474629,-474626,-474623,-474620,-474616,-474613,-474610,-474607,-474604,-474601,-474598,-474595,-474592,-474589,-474585,-474582,-474579,-474576,-474573,-474570,-474567,-474564,-474561,-474557,-474554,-474551,-474548,-474545,-474542,-474539,-474536,-474533,-474530,-474526,-474523,-474520,-474517,-474514,-474511,-474508,-474505,-474502,-474498,-474495,-474492,-474489,-474486,-474483,-474480,-474477,-474474,-474471,-474467,-474464,-474461,-474458,-474455,-474452,-474449,-474446,-474443,-474439,-474436,-474433,-474430,-474427,-474424,-474421,-474418,-474415,-474411,-474408,-474405,-474402,-474399,-474396,-474393,-474390,-474387,-474383,-474380,-474377,-474374,-474371,-474368,-474365,-474362,-474359,-474355,-474352,-474349,-474346,-474343,-474340,-474337,-474334,-474331,-474327,-474324,-474321,-474318,-474315,-474312,-474309,-474306,-474302,-474299,-474296,-474293,-474290,-474287,-474284,-474281,-474278,-474274,-474271,-474268,-474265,-474262,-474259,-474256,-474253,-474250,-474246,-474243,-474240,-474237,-474234,-474231,-474228,-474225,-474221,-474218,-474215,-474212,-474209,-474206,-474203,-474200,-474196,-474193,-474190,-474187,-474184,-474181,-474178,-474175,-474172,-474168,-474165,-474162,-474159,-474156,-474153,-474150,-474147,-474143,-474140,-474137,-474134,-474131,-474128,-474125,-474122,-474118,-474115,-474112,-474109,-474106,-474103,-474100,-474097,-474093,-474090,-474087,-474084,-474081,-474078,-474075,-474072,-474068,-474065,-474062,-474059,-474056,-474053,-474050,-474047,-474043,-474040,-474037,-474034,-474031,-474028,-474025,-474022,-474018,-474015,-474012,-474009,-474006,-474003,-474000,-473997,-473993,-473990,-473987,-473984,-473981,-473978,-473975,-473972,-473968,-473965,-473962,-473959,-473956,-473953,-473950,-473947,-473943,-473940,-473937,-473934,-473931,-473928,-473925,-473921,-473918,-473915,-473912,-473909,-473906,-473903,-473900,-473896,-473893,-473890,-473887,-473884,-473881,-473878,-473875,-473871,-473868,-473865,-473862,-473859,-473856,-473853,-473849,-473846,-473843,-473840,-473837,-473834,-473831,-473828,-473824,-473821,-473818,-473815,-473812,-473809,-473806,-473802,-473799,-473796,-473793,-473790,-473787,-473784,-473780,-473777,-473774,-473771,-473768,-473765,-473762,-473759,-473755,-473752,-473749,-473746,-473743,-473740,-473737,-473733,-473730,-473727,-473724,-473721,-473718,-473715,-473711,-473708,-473705,-473702,-473699,-473696,-473693,-473689,-473686,-473683,-473680,-473677,-473674,-473671,-473668,-473664,-473661,-473658,-473655,-473652,-473649,-473646,-473642,-473639,-473636,-473633,-473630,-473627,-473624,-473620,-473617,-473614,-473611,-473608,-473605,-473602,-473598,-473595,-473592,-473589,-473586,-473583,-473580,-473576,-473573,-473570,-473567,-473564,-473561,-473557,-473554,-473551,-473548,-473545,-473542,-473539,-473535,-473532,-473529,-473526,-473523,-473520,-473517,-473513,-473510,-473507,-473504,-473501,-473498,-473495,-473491,-473488,-473485,-473482,-473479,-473476,-473473,-473469,-473466,-473463,-473460,-473457,-473454,-473450,-473447,-473444,-473441,-473438,-473435,-473432,-473428,-473425,-473422,-473419,-473416,-473413,-473410,-473406,-473403,-473400,-473397,-473394,-473391,-473387,-473384,-473381,-473378,-473375,-473372,-473369,-473365,-473362,-473359,-473356,-473353,-473350,-473346,-473343,-473340,-473337,-473334,-473331,-473328,-473324,-473321,-473318,-473315,-473312,-473309,-473305,-473302,-473299,-473296,-473293,-473290,-473287,-473283,-473280,-473277,-473274,-473271,-473268,-473264,-473261,-473258,-473255,-473252,-473249,-473245,-473242,-473239,-473236,-473233,-473230,-473227,-473223,-473220,-473217,-473214,-473211,-473208,-473204,-473201,-473198,-473195,-473192,-473189,-473185,-473182,-473179,-473176,-473173,-473170,-473167,-473163,-473160,-473157,-473154,-473151,-473148,-473144,-473141,-473138,-473135,-473132,-473129,-473125,-473122,-473119,-473116,-473113,-473110,-473106,-473103,-473100,-473097,-473094,-473091,-473087,-473084,-473081,-473078,-473075,-473072,-473068,-473065,-473062,-473059,-473056,-473053,-473049,-473046,-473043,-473040,-473037,-473034,-473030,-473027,-473024,-473021,-473018,-473015,-473011,-473008,-473005,-473002,-472999,-472996,-472992,-472989,-472986,-472983,-472980,-472977,-472973,-472970,-472967,-472964,-472961,-472958,-472954,-472951,-472948,-472945,-472942,-472939,-472935,-472932,-472929,-472926,-472923,-472920,-472916,-472913,-472910,-472907,-472904,-472901,-472897,-472894,-472891,-472888,-472885,-472882,-472878,-472875,-472872,-472869,-472866,-472862,-472859,-472856,-472853,-472850,-472847,-472843,-472840,-472837,-472834,-472831,-472828,-472824,-472821,-472818,-472815,-472812,-472809,-472805,-472802,-472799,-472796,-472793,-472789,-472786,-472783,-472780,-472777,-472774,-472770,-472767,-472764,-472761,-472758,-472755,-472751,-472748,-472745,-472742,-472739,-472735,-472732,-472729,-472726,-472723,-472720,-472716,-472713,-472710,-472707,-472704,-472700,-472697,-472694,-472691,-472688,-472685,-472681,-472678,-472675,-472672,-472669,-472665,-472662,-472659,-472656,-472653,-472650,-472646,-472643,-472640,-472637,-472634,-472630,-472627,-472624,-472621,-472618,-472615,-472611,-472608,-472605,-472602,-472599,-472595,-472592,-472589,-472586,-472583,-472580,-472576,-472573,-472570,-472567,-472564,-472560,-472557,-472554,-472551,-472548,-472545,-472541,-472538,-472535,-472532,-472529,-472525,-472522,-472519,-472516,-472513,-472509,-472506,-472503,-472500,-472497,-472494,-472490,-472487,-472484,-472481,-472478,-472474,-472471,-472468,-472465,-472462,-472458,-472455,-472452,-472449,-472446,-472443,-472439,-472436,-472433,-472430,-472427,-472423,-472420,-472417,-472414,-472411,-472407,-472404,-472401,-472398,-472395,-472391,-472388,-472385,-472382,-472379,-472375,-472372,-472369,-472366,-472363,-472360,-472356,-472353,-472350,-472347,-472344,-472340,-472337,-472334,-472331,-472328,-472324,-472321,-472318,-472315,-472312,-472308,-472305,-472302,-472299,-472296,-472292,-472289,-472286,-472283,-472280,-472276,-472273,-472270,-472267,-472264,-472260,-472257,-472254,-472251,-472248,-472244,-472241,-472238,-472235,-472232,-472229,-472225,-472222,-472219,-472216,-472213,-472209,-472206,-472203,-472200,-472197,-472193,-472190,-472187,-472184,-472181,-472177 
);

type cA2_array_type is array (0 to Arr_size) of integer;
signal A2 : cA2_array_type:= (others => 248765);

type cB0_array_type is array (0 to Arr_size) of integer;
signal B0 : cB0_array_type:= (others =>248765);

type cB1_array_type is array (0 to Arr_size) of integer;
signal B1 : cB1_array_type:= (others => 6689);

type cB2_array_type is array (0 to Arr_size) of integer;
signal B2 : cB2_array_type:=(others => -6689);

signal constA0 : signed(w_coef-1 downto 0):= to_signed(A0(0),w_coef);
signal constA1 : signed(w_coef-1 downto 0):= to_signed(A1(0),w_coef);
signal constA2 : signed(w_coef-1 downto 0):= to_signed(A2(0),w_coef);
signal constB0 : signed(w_coef-1 downto 0) := to_signed(B0(0),w_coef);
signal constB1 : signed(w_coef-1 downto 0):= to_signed(B1(0),w_coef);
signal constB2 : signed(w_coef-1 downto 0):= to_signed(B2(0),w_coef);

signal BP_out : signed(W_in-1 downto 0) := (others =>'0');
signal data_out_temp:  signed(W_in-1 downto 0) := (others =>'0');
signal BW_clk : std_logic := '0';
begin

process(CLK_50,nReset) 
variable counter : integer := 0;
variable direction: std_logic := '0';
begin
if (nReset = '0') then
	counter := 0;
	direction:= '0';
elsif (rising_edge(CLK_50)) then
	data_out_temp <= BP_out+data_in; -- output 
	if (new_val = '1') then
	if (direction = '0') then
		constA0 <= to_signed(A0(counter),w_coef);
		constA1 <= to_signed(A1(counter),w_coef);
		constA2 <= to_signed(A2(counter),w_coef);
		constB0 <= to_signed(B0(counter),w_coef);
		constB1 <= to_signed(B1(counter),w_coef);
		constB2 <= to_signed(B2(counter),w_coef);
		counter := counter + 1;
		if(counter = Arr_size) then
			direction := '1';
		end if;
	end if;
	if(direction = '1') then
		counter := counter -1;
		constA0 <= to_signed(A0(counter),w_coef);
		constA1 <= to_signed(A1(counter),w_coef);
		constA2 <= to_signed(A2(counter),w_coef);
		constB0 <= to_signed(B0(counter),w_coef);
		constB1 <= to_signed(B1(counter),w_coef);
		constB2 <= to_signed(B2(counter),w_coef);
		if(counter = 0) then
			direction := '0';
		end if;
	end if;
	end if;
end if;
end process;

IIRDF_inst : IIRDF1_BW 
generic map(
    W_in => W_in,
	 W_coef => W_coef

)
port map(
	iCLK => CLK_50,          
	iRESET_N => nReset,      
	new_val => new_val,        
	IIR_in => data_in,                 
	IIR_out => BP_out ,        

	B0 => constB0,
   B1 => constB1,
   B2 => constB2,
   A0 => constA0,
   A1 => constA1,
   A2 => constA2
);

process(CLK_50,nReset)
begin
if nReset = '0' then
	data_out <= (others => '0');
elsif(rising_edge(CLK_50)) then
	if(new_val = '1') then
	if WahWah_EN = '0' then
		data_out <= data_in;
	elsif WahWah_EN = '1' then
		data_out <= shift_right(data_out_temp + data_in,1);
	end if;
	end if;
end if;
end process;
end;