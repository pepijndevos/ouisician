library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity WahWah_FX is
port (
	CLK_50		: in std_logic;
	nReset		: in std_logic;
	new_val		: in std_logic;       -- indicates a new input value, input from data_over
	data_in		: in signed (15 downto 0);         
	data_out		: out signed (15 downto 0);   -- Output
	WahWah_EN 	: in std_logic
);
end entity WahWah_FX;

architecture behaviour of WahWah_FX is
constant W_coef : integer := 23;
constant W_in : integer := 16;
constant A0 : integer :=1048576 ;
constant A2 : integer :=1034939 ;
constant B0 : integer :=6818 ;
constant B1 : integer := 0;
constant B2 : integer := -6818 ; 
constant Arr_size : integer := 24000;

component IIRDF1_BW is
generic (
   W_in : integer ;
	W_coef : integer;
	A0 : integer;
	A2 : integer;
	B0 : integer ;
	B1 : integer;
	B2 : integer    
);
port (
	iCLK            : in std_logic;
	iRESET_N        : in std_logic;
	new_val         : in std_logic;       -- indicates a new input value, input from data_over
	IIR_in          : in signed (15 downto 0);   -- singed is expected             
	IIR_out         : out signed (15 downto 0);   -- Output
   A1 : in signed(W_coef-1 downto 0)

);
end component;


type cA1_array_type is array (0 to Arr_size) of integer;
signal A1 : cA1_array_type:=(-2079097,-2079095,-2079093,-2079091,-2079089,-2079088,-2079086,-2079084,-2079082,-2079080,-2079078,-2079076,-2079075,-2079073,-2079071,-2079069,-2079067,-2079065,-2079063,-2079062,-2079060,-2079058,-2079056,-2079054,-2079052,-2079050,-2079048,-2079047,-2079045,-2079043,-2079041,-2079039,-2079037,-2079035,-2079034,-2079032,-2079030,-2079028,-2079026,-2079024,-2079022,-2079020,-2079019,-2079017,-2079015,-2079013,-2079011,-2079009,-2079007,-2079005,-2079004,-2079002,-2079000,-2078998,-2078996,-2078994,-2078992,-2078990,-2078988,-2078987,-2078985,-2078983,-2078981,-2078979,-2078977,-2078975,-2078973,-2078972,-2078970,-2078968,-2078966,-2078964,-2078962,-2078960,-2078958,-2078956,-2078955,-2078953,-2078951,-2078949,-2078947,-2078945,-2078943,-2078941,-2078939,-2078938,-2078936,-2078934,-2078932,-2078930,-2078928,-2078926,-2078924,-2078922,-2078921,-2078919,-2078917,-2078915,-2078913,-2078911,-2078909,-2078907,-2078905,-2078903,-2078902,-2078900,-2078898,-2078896,-2078894,-2078892,-2078890,-2078888,-2078886,-2078884,-2078883,-2078881,-2078879,-2078877,-2078875,-2078873,-2078871,-2078869,-2078867,-2078865,-2078864,-2078862,-2078860,-2078858,-2078856,-2078854,-2078852,-2078850,-2078848,-2078846,-2078844,-2078843,-2078841,-2078839,-2078837,-2078835,-2078833,-2078831,-2078829,-2078827,-2078825,-2078823,-2078821,-2078820,-2078818,-2078816,-2078814,-2078812,-2078810,-2078808,-2078806,-2078804,-2078802,-2078800,-2078798,-2078797,-2078795,-2078793,-2078791,-2078789,-2078787,-2078785,-2078783,-2078781,-2078779,-2078777,-2078775,-2078773,-2078772,-2078770,-2078768,-2078766,-2078764,-2078762,-2078760,-2078758,-2078756,-2078754,-2078752,-2078750,-2078748,-2078746,-2078745,-2078743,-2078741,-2078739,-2078737,-2078735,-2078733,-2078731,-2078729,-2078727,-2078725,-2078723,-2078721,-2078719,-2078718,-2078716,-2078714,-2078712,-2078710,-2078708,-2078706,-2078704,-2078702,-2078700,-2078698,-2078696,-2078694,-2078692,-2078690,-2078688,-2078686,-2078685,-2078683,-2078681,-2078679,-2078677,-2078675,-2078673,-2078671,-2078669,-2078667,-2078665,-2078663,-2078661,-2078659,-2078657,-2078655,-2078653,-2078651,-2078650,-2078648,-2078646,-2078644,-2078642,-2078640,-2078638,-2078636,-2078634,-2078632,-2078630,-2078628,-2078626,-2078624,-2078622,-2078620,-2078618,-2078616,-2078614,-2078612,-2078610,-2078608,-2078607,-2078605,-2078603,-2078601,-2078599,-2078597,-2078595,-2078593,-2078591,-2078589,-2078587,-2078585,-2078583,-2078581,-2078579,-2078577,-2078575,-2078573,-2078571,-2078569,-2078567,-2078565,-2078563,-2078561,-2078559,-2078557,-2078556,-2078554,-2078552,-2078550,-2078548,-2078546,-2078544,-2078542,-2078540,-2078538,-2078536,-2078534,-2078532,-2078530,-2078528,-2078526,-2078524,-2078522,-2078520,-2078518,-2078516,-2078514,-2078512,-2078510,-2078508,-2078506,-2078504,-2078502,-2078500,-2078498,-2078496,-2078494,-2078492,-2078490,-2078488,-2078486,-2078484,-2078482,-2078480,-2078478,-2078476,-2078474,-2078473,-2078471,-2078469,-2078467,-2078465,-2078463,-2078461,-2078459,-2078457,-2078455,-2078453,-2078451,-2078449,-2078447,-2078445,-2078443,-2078441,-2078439,-2078437,-2078435,-2078433,-2078431,-2078429,-2078427,-2078425,-2078423,-2078421,-2078419,-2078417,-2078415,-2078413,-2078411,-2078409,-2078407,-2078405,-2078403,-2078401,-2078399,-2078397,-2078395,-2078393,-2078391,-2078389,-2078387,-2078385,-2078383,-2078381,-2078379,-2078377,-2078375,-2078373,-2078371,-2078369,-2078367,-2078365,-2078363,-2078361,-2078359,-2078357,-2078355,-2078353,-2078351,-2078349,-2078347,-2078345,-2078343,-2078341,-2078339,-2078337,-2078335,-2078333,-2078331,-2078329,-2078327,-2078325,-2078323,-2078321,-2078319,-2078317,-2078315,-2078313,-2078311,-2078309,-2078306,-2078304,-2078302,-2078300,-2078298,-2078296,-2078294,-2078292,-2078290,-2078288,-2078286,-2078284,-2078282,-2078280,-2078278,-2078276,-2078274,-2078272,-2078270,-2078268,-2078266,-2078264,-2078262,-2078260,-2078258,-2078256,-2078254,-2078252,-2078250,-2078248,-2078246,-2078244,-2078242,-2078240,-2078238,-2078236,-2078234,-2078232,-2078230,-2078228,-2078226,-2078224,-2078221,-2078219,-2078217,-2078215,-2078213,-2078211,-2078209,-2078207,-2078205,-2078203,-2078201,-2078199,-2078197,-2078195,-2078193,-2078191,-2078189,-2078187,-2078185,-2078183,-2078181,-2078179,-2078177,-2078175,-2078173,-2078171,-2078169,-2078166,-2078164,-2078162,-2078160,-2078158,-2078156,-2078154,-2078152,-2078150,-2078148,-2078146,-2078144,-2078142,-2078140,-2078138,-2078136,-2078134,-2078132,-2078130,-2078128,-2078126,-2078123,-2078121,-2078119,-2078117,-2078115,-2078113,-2078111,-2078109,-2078107,-2078105,-2078103,-2078101,-2078099,-2078097,-2078095,-2078093,-2078091,-2078089,-2078086,-2078084,-2078082,-2078080,-2078078,-2078076,-2078074,-2078072,-2078070,-2078068,-2078066,-2078064,-2078062,-2078060,-2078058,-2078056,-2078054,-2078051,-2078049,-2078047,-2078045,-2078043,-2078041,-2078039,-2078037,-2078035,-2078033,-2078031,-2078029,-2078027,-2078025,-2078023,-2078020,-2078018,-2078016,-2078014,-2078012,-2078010,-2078008,-2078006,-2078004,-2078002,-2078000,-2077998,-2077996,-2077994,-2077991,-2077989,-2077987,-2077985,-2077983,-2077981,-2077979,-2077977,-2077975,-2077973,-2077971,-2077969,-2077966,-2077964,-2077962,-2077960,-2077958,-2077956,-2077954,-2077952,-2077950,-2077948,-2077946,-2077944,-2077941,-2077939,-2077937,-2077935,-2077933,-2077931,-2077929,-2077927,-2077925,-2077923,-2077921,-2077919,-2077916,-2077914,-2077912,-2077910,-2077908,-2077906,-2077904,-2077902,-2077900,-2077898,-2077896,-2077893,-2077891,-2077889,-2077887,-2077885,-2077883,-2077881,-2077879,-2077877,-2077875,-2077872,-2077870,-2077868,-2077866,-2077864,-2077862,-2077860,-2077858,-2077856,-2077854,-2077851,-2077849,-2077847,-2077845,-2077843,-2077841,-2077839,-2077837,-2077835,-2077833,-2077830,-2077828,-2077826,-2077824,-2077822,-2077820,-2077818,-2077816,-2077814,-2077811,-2077809,-2077807,-2077805,-2077803,-2077801,-2077799,-2077797,-2077795,-2077792,-2077790,-2077788,-2077786,-2077784,-2077782,-2077780,-2077778,-2077776,-2077773,-2077771,-2077769,-2077767,-2077765,-2077763,-2077761,-2077759,-2077757,-2077754,-2077752,-2077750,-2077748,-2077746,-2077744,-2077742,-2077740,-2077737,-2077735,-2077733,-2077731,-2077729,-2077727,-2077725,-2077723,-2077720,-2077718,-2077716,-2077714,-2077712,-2077710,-2077708,-2077706,-2077703,-2077701,-2077699,-2077697,-2077695,-2077693,-2077691,-2077689,-2077686,-2077684,-2077682,-2077680,-2077678,-2077676,-2077674,-2077671,-2077669,-2077667,-2077665,-2077663,-2077661,-2077659,-2077657,-2077654,-2077652,-2077650,-2077648,-2077646,-2077644,-2077642,-2077639,-2077637,-2077635,-2077633,-2077631,-2077629,-2077627,-2077624,-2077622,-2077620,-2077618,-2077616,-2077614,-2077612,-2077609,-2077607,-2077605,-2077603,-2077601,-2077599,-2077597,-2077594,-2077592,-2077590,-2077588,-2077586,-2077584,-2077581,-2077579,-2077577,-2077575,-2077573,-2077571,-2077569,-2077566,-2077564,-2077562,-2077560,-2077558,-2077556,-2077553,-2077551,-2077549,-2077547,-2077545,-2077543,-2077541,-2077538,-2077536,-2077534,-2077532,-2077530,-2077528,-2077525,-2077523,-2077521,-2077519,-2077517,-2077515,-2077512,-2077510,-2077508,-2077506,-2077504,-2077502,-2077499,-2077497,-2077495,-2077493,-2077491,-2077489,-2077486,-2077484,-2077482,-2077480,-2077478,-2077476,-2077473,-2077471,-2077469,-2077467,-2077465,-2077463,-2077460,-2077458,-2077456,-2077454,-2077452,-2077450,-2077447,-2077445,-2077443,-2077441,-2077439,-2077437,-2077434,-2077432,-2077430,-2077428,-2077426,-2077423,-2077421,-2077419,-2077417,-2077415,-2077413,-2077410,-2077408,-2077406,-2077404,-2077402,-2077399,-2077397,-2077395,-2077393,-2077391,-2077389,-2077386,-2077384,-2077382,-2077380,-2077378,-2077375,-2077373,-2077371,-2077369,-2077367,-2077364,-2077362,-2077360,-2077358,-2077356,-2077354,-2077351,-2077349,-2077347,-2077345,-2077343,-2077340,-2077338,-2077336,-2077334,-2077332,-2077329,-2077327,-2077325,-2077323,-2077321,-2077318,-2077316,-2077314,-2077312,-2077310,-2077307,-2077305,-2077303,-2077301,-2077299,-2077296,-2077294,-2077292,-2077290,-2077288,-2077285,-2077283,-2077281,-2077279,-2077277,-2077274,-2077272,-2077270,-2077268,-2077266,-2077263,-2077261,-2077259,-2077257,-2077255,-2077252,-2077250,-2077248,-2077246,-2077243,-2077241,-2077239,-2077237,-2077235,-2077232,-2077230,-2077228,-2077226,-2077224,-2077221,-2077219,-2077217,-2077215,-2077213,-2077210,-2077208,-2077206,-2077204,-2077201,-2077199,-2077197,-2077195,-2077193,-2077190,-2077188,-2077186,-2077184,-2077181,-2077179,-2077177,-2077175,-2077173,-2077170,-2077168,-2077166,-2077164,-2077161,-2077159,-2077157,-2077155,-2077153,-2077150,-2077148,-2077146,-2077144,-2077141,-2077139,-2077137,-2077135,-2077132,-2077130,-2077128,-2077126,-2077124,-2077121,-2077119,-2077117,-2077115,-2077112,-2077110,-2077108,-2077106,-2077103,-2077101,-2077099,-2077097,-2077095,-2077092,-2077090,-2077088,-2077086,-2077083,-2077081,-2077079,-2077077,-2077074,-2077072,-2077070,-2077068,-2077065,-2077063,-2077061,-2077059,-2077056,-2077054,-2077052,-2077050,-2077047,-2077045,-2077043,-2077041,-2077038,-2077036,-2077034,-2077032,-2077029,-2077027,-2077025,-2077023,-2077021,-2077018,-2077016,-2077014,-2077012,-2077009,-2077007,-2077005,-2077002,-2077000,-2076998,-2076996,-2076993,-2076991,-2076989,-2076987,-2076984,-2076982,-2076980,-2076978,-2076975,-2076973,-2076971,-2076969,-2076966,-2076964,-2076962,-2076960,-2076957,-2076955,-2076953,-2076951,-2076948,-2076946,-2076944,-2076942,-2076939,-2076937,-2076935,-2076932,-2076930,-2076928,-2076926,-2076923,-2076921,-2076919,-2076917,-2076914,-2076912,-2076910,-2076908,-2076905,-2076903,-2076901,-2076898,-2076896,-2076894,-2076892,-2076889,-2076887,-2076885,-2076883,-2076880,-2076878,-2076876,-2076873,-2076871,-2076869,-2076867,-2076864,-2076862,-2076860,-2076858,-2076855,-2076853,-2076851,-2076848,-2076846,-2076844,-2076842,-2076839,-2076837,-2076835,-2076832,-2076830,-2076828,-2076826,-2076823,-2076821,-2076819,-2076817,-2076814,-2076812,-2076810,-2076807,-2076805,-2076803,-2076801,-2076798,-2076796,-2076794,-2076791,-2076789,-2076787,-2076785,-2076782,-2076780,-2076778,-2076775,-2076773,-2076771,-2076768,-2076766,-2076764,-2076762,-2076759,-2076757,-2076755,-2076752,-2076750,-2076748,-2076746,-2076743,-2076741,-2076739,-2076736,-2076734,-2076732,-2076729,-2076727,-2076725,-2076723,-2076720,-2076718,-2076716,-2076713,-2076711,-2076709,-2076706,-2076704,-2076702,-2076700,-2076697,-2076695,-2076693,-2076690,-2076688,-2076686,-2076683,-2076681,-2076679,-2076676,-2076674,-2076672,-2076670,-2076667,-2076665,-2076663,-2076660,-2076658,-2076656,-2076653,-2076651,-2076649,-2076646,-2076644,-2076642,-2076640,-2076637,-2076635,-2076633,-2076630,-2076628,-2076626,-2076623,-2076621,-2076619,-2076616,-2076614,-2076612,-2076609,-2076607,-2076605,-2076602,-2076600,-2076598,-2076595,-2076593,-2076591,-2076589,-2076586,-2076584,-2076582,-2076579,-2076577,-2076575,-2076572,-2076570,-2076568,-2076565,-2076563,-2076561,-2076558,-2076556,-2076554,-2076551,-2076549,-2076547,-2076544,-2076542,-2076540,-2076537,-2076535,-2076533,-2076530,-2076528,-2076526,-2076523,-2076521,-2076519,-2076516,-2076514,-2076512,-2076509,-2076507,-2076505,-2076502,-2076500,-2076498,-2076495,-2076493,-2076491,-2076488,-2076486,-2076484,-2076481,-2076479,-2076477,-2076474,-2076472,-2076470,-2076467,-2076465,-2076463,-2076460,-2076458,-2076456,-2076453,-2076451,-2076449,-2076446,-2076444,-2076441,-2076439,-2076437,-2076434,-2076432,-2076430,-2076427,-2076425,-2076423,-2076420,-2076418,-2076416,-2076413,-2076411,-2076409,-2076406,-2076404,-2076402,-2076399,-2076397,-2076394,-2076392,-2076390,-2076387,-2076385,-2076383,-2076380,-2076378,-2076376,-2076373,-2076371,-2076369,-2076366,-2076364,-2076361,-2076359,-2076357,-2076354,-2076352,-2076350,-2076347,-2076345,-2076343,-2076340,-2076338,-2076335,-2076333,-2076331,-2076328,-2076326,-2076324,-2076321,-2076319,-2076317,-2076314,-2076312,-2076309,-2076307,-2076305,-2076302,-2076300,-2076298,-2076295,-2076293,-2076291,-2076288,-2076286,-2076283,-2076281,-2076279,-2076276,-2076274,-2076272,-2076269,-2076267,-2076264,-2076262,-2076260,-2076257,-2076255,-2076253,-2076250,-2076248,-2076245,-2076243,-2076241,-2076238,-2076236,-2076233,-2076231,-2076229,-2076226,-2076224,-2076222,-2076219,-2076217,-2076214,-2076212,-2076210,-2076207,-2076205,-2076203,-2076200,-2076198,-2076195,-2076193,-2076191,-2076188,-2076186,-2076183,-2076181,-2076179,-2076176,-2076174,-2076171,-2076169,-2076167,-2076164,-2076162,-2076160,-2076157,-2076155,-2076152,-2076150,-2076148,-2076145,-2076143,-2076140,-2076138,-2076136,-2076133,-2076131,-2076128,-2076126,-2076124,-2076121,-2076119,-2076116,-2076114,-2076112,-2076109,-2076107,-2076104,-2076102,-2076100,-2076097,-2076095,-2076092,-2076090,-2076088,-2076085,-2076083,-2076080,-2076078,-2076076,-2076073,-2076071,-2076068,-2076066,-2076064,-2076061,-2076059,-2076056,-2076054,-2076051,-2076049,-2076047,-2076044,-2076042,-2076039,-2076037,-2076035,-2076032,-2076030,-2076027,-2076025,-2076023,-2076020,-2076018,-2076015,-2076013,-2076010,-2076008,-2076006,-2076003,-2076001,-2075998,-2075996,-2075994,-2075991,-2075989,-2075986,-2075984,-2075981,-2075979,-2075977,-2075974,-2075972,-2075969,-2075967,-2075964,-2075962,-2075960,-2075957,-2075955,-2075952,-2075950,-2075947,-2075945,-2075943,-2075940,-2075938,-2075935,-2075933,-2075930,-2075928,-2075926,-2075923,-2075921,-2075918,-2075916,-2075913,-2075911,-2075909,-2075906,-2075904,-2075901,-2075899,-2075896,-2075894,-2075892,-2075889,-2075887,-2075884,-2075882,-2075879,-2075877,-2075875,-2075872,-2075870,-2075867,-2075865,-2075862,-2075860,-2075857,-2075855,-2075853,-2075850,-2075848,-2075845,-2075843,-2075840,-2075838,-2075835,-2075833,-2075831,-2075828,-2075826,-2075823,-2075821,-2075818,-2075816,-2075813,-2075811,-2075809,-2075806,-2075804,-2075801,-2075799,-2075796,-2075794,-2075791,-2075789,-2075787,-2075784,-2075782,-2075779,-2075777,-2075774,-2075772,-2075769,-2075767,-2075764,-2075762,-2075760,-2075757,-2075755,-2075752,-2075750,-2075747,-2075745,-2075742,-2075740,-2075737,-2075735,-2075732,-2075730,-2075728,-2075725,-2075723,-2075720,-2075718,-2075715,-2075713,-2075710,-2075708,-2075705,-2075703,-2075700,-2075698,-2075696,-2075693,-2075691,-2075688,-2075686,-2075683,-2075681,-2075678,-2075676,-2075673,-2075671,-2075668,-2075666,-2075663,-2075661,-2075658,-2075656,-2075654,-2075651,-2075649,-2075646,-2075644,-2075641,-2075639,-2075636,-2075634,-2075631,-2075629,-2075626,-2075624,-2075621,-2075619,-2075616,-2075614,-2075611,-2075609,-2075607,-2075604,-2075602,-2075599,-2075597,-2075594,-2075592,-2075589,-2075587,-2075584,-2075582,-2075579,-2075577,-2075574,-2075572,-2075569,-2075567,-2075564,-2075562,-2075559,-2075557,-2075554,-2075552,-2075549,-2075547,-2075544,-2075542,-2075539,-2075537,-2075534,-2075532,-2075529,-2075527,-2075524,-2075522,-2075519,-2075517,-2075514,-2075512,-2075509,-2075507,-2075504,-2075502,-2075500,-2075497,-2075495,-2075492,-2075490,-2075487,-2075485,-2075482,-2075480,-2075477,-2075475,-2075472,-2075470,-2075467,-2075465,-2075462,-2075460,-2075457,-2075455,-2075452,-2075449,-2075447,-2075444,-2075442,-2075439,-2075437,-2075434,-2075432,-2075429,-2075427,-2075424,-2075422,-2075419,-2075417,-2075414,-2075412,-2075409,-2075407,-2075404,-2075402,-2075399,-2075397,-2075394,-2075392,-2075389,-2075387,-2075384,-2075382,-2075379,-2075377,-2075374,-2075372,-2075369,-2075367,-2075364,-2075362,-2075359,-2075357,-2075354,-2075352,-2075349,-2075346,-2075344,-2075341,-2075339,-2075336,-2075334,-2075331,-2075329,-2075326,-2075324,-2075321,-2075319,-2075316,-2075314,-2075311,-2075309,-2075306,-2075304,-2075301,-2075299,-2075296,-2075293,-2075291,-2075288,-2075286,-2075283,-2075281,-2075278,-2075276,-2075273,-2075271,-2075268,-2075266,-2075263,-2075261,-2075258,-2075256,-2075253,-2075250,-2075248,-2075245,-2075243,-2075240,-2075238,-2075235,-2075233,-2075230,-2075228,-2075225,-2075223,-2075220,-2075217,-2075215,-2075212,-2075210,-2075207,-2075205,-2075202,-2075200,-2075197,-2075195,-2075192,-2075190,-2075187,-2075184,-2075182,-2075179,-2075177,-2075174,-2075172,-2075169,-2075167,-2075164,-2075162,-2075159,-2075156,-2075154,-2075151,-2075149,-2075146,-2075144,-2075141,-2075139,-2075136,-2075133,-2075131,-2075128,-2075126,-2075123,-2075121,-2075118,-2075116,-2075113,-2075110,-2075108,-2075105,-2075103,-2075100,-2075098,-2075095,-2075093,-2075090,-2075087,-2075085,-2075082,-2075080,-2075077,-2075075,-2075072,-2075070,-2075067,-2075064,-2075062,-2075059,-2075057,-2075054,-2075052,-2075049,-2075046,-2075044,-2075041,-2075039,-2075036,-2075034,-2075031,-2075028,-2075026,-2075023,-2075021,-2075018,-2075016,-2075013,-2075010,-2075008,-2075005,-2075003,-2075000,-2074998,-2074995,-2074992,-2074990,-2074987,-2074985,-2074982,-2074980,-2074977,-2074974,-2074972,-2074969,-2074967,-2074964,-2074962,-2074959,-2074956,-2074954,-2074951,-2074949,-2074946,-2074944,-2074941,-2074938,-2074936,-2074933,-2074931,-2074928,-2074925,-2074923,-2074920,-2074918,-2074915,-2074913,-2074910,-2074907,-2074905,-2074902,-2074900,-2074897,-2074894,-2074892,-2074889,-2074887,-2074884,-2074881,-2074879,-2074876,-2074874,-2074871,-2074868,-2074866,-2074863,-2074861,-2074858,-2074856,-2074853,-2074850,-2074848,-2074845,-2074843,-2074840,-2074837,-2074835,-2074832,-2074830,-2074827,-2074824,-2074822,-2074819,-2074817,-2074814,-2074811,-2074809,-2074806,-2074804,-2074801,-2074798,-2074796,-2074793,-2074791,-2074788,-2074785,-2074783,-2074780,-2074778,-2074775,-2074772,-2074770,-2074767,-2074764,-2074762,-2074759,-2074757,-2074754,-2074751,-2074749,-2074746,-2074744,-2074741,-2074738,-2074736,-2074733,-2074731,-2074728,-2074725,-2074723,-2074720,-2074717,-2074715,-2074712,-2074710,-2074707,-2074704,-2074702,-2074699,-2074697,-2074694,-2074691,-2074689,-2074686,-2074683,-2074681,-2074678,-2074676,-2074673,-2074670,-2074668,-2074665,-2074663,-2074660,-2074657,-2074655,-2074652,-2074649,-2074647,-2074644,-2074642,-2074639,-2074636,-2074634,-2074631,-2074628,-2074626,-2074623,-2074620,-2074618,-2074615,-2074613,-2074610,-2074607,-2074605,-2074602,-2074599,-2074597,-2074594,-2074592,-2074589,-2074586,-2074584,-2074581,-2074578,-2074576,-2074573,-2074570,-2074568,-2074565,-2074563,-2074560,-2074557,-2074555,-2074552,-2074549,-2074547,-2074544,-2074541,-2074539,-2074536,-2074534,-2074531,-2074528,-2074526,-2074523,-2074520,-2074518,-2074515,-2074512,-2074510,-2074507,-2074504,-2074502,-2074499,-2074497,-2074494,-2074491,-2074489,-2074486,-2074483,-2074481,-2074478,-2074475,-2074473,-2074470,-2074467,-2074465,-2074462,-2074459,-2074457,-2074454,-2074451,-2074449,-2074446,-2074443,-2074441,-2074438,-2074436,-2074433,-2074430,-2074428,-2074425,-2074422,-2074420,-2074417,-2074414,-2074412,-2074409,-2074406,-2074404,-2074401,-2074398,-2074396,-2074393,-2074390,-2074388,-2074385,-2074382,-2074380,-2074377,-2074374,-2074372,-2074369,-2074366,-2074364,-2074361,-2074358,-2074356,-2074353,-2074350,-2074348,-2074345,-2074342,-2074340,-2074337,-2074334,-2074332,-2074329,-2074326,-2074324,-2074321,-2074318,-2074316,-2074313,-2074310,-2074308,-2074305,-2074302,-2074300,-2074297,-2074294,-2074292,-2074289,-2074286,-2074284,-2074281,-2074278,-2074275,-2074273,-2074270,-2074267,-2074265,-2074262,-2074259,-2074257,-2074254,-2074251,-2074249,-2074246,-2074243,-2074241,-2074238,-2074235,-2074233,-2074230,-2074227,-2074225,-2074222,-2074219,-2074216,-2074214,-2074211,-2074208,-2074206,-2074203,-2074200,-2074198,-2074195,-2074192,-2074190,-2074187,-2074184,-2074181,-2074179,-2074176,-2074173,-2074171,-2074168,-2074165,-2074163,-2074160,-2074157,-2074155,-2074152,-2074149,-2074146,-2074144,-2074141,-2074138,-2074136,-2074133,-2074130,-2074128,-2074125,-2074122,-2074119,-2074117,-2074114,-2074111,-2074109,-2074106,-2074103,-2074101,-2074098,-2074095,-2074092,-2074090,-2074087,-2074084,-2074082,-2074079,-2074076,-2074073,-2074071,-2074068,-2074065,-2074063,-2074060,-2074057,-2074054,-2074052,-2074049,-2074046,-2074044,-2074041,-2074038,-2074036,-2074033,-2074030,-2074027,-2074025,-2074022,-2074019,-2074017,-2074014,-2074011,-2074008,-2074006,-2074003,-2074000,-2073997,-2073995,-2073992,-2073989,-2073987,-2073984,-2073981,-2073978,-2073976,-2073973,-2073970,-2073968,-2073965,-2073962,-2073959,-2073957,-2073954,-2073951,-2073948,-2073946,-2073943,-2073940,-2073938,-2073935,-2073932,-2073929,-2073927,-2073924,-2073921,-2073918,-2073916,-2073913,-2073910,-2073908,-2073905,-2073902,-2073899,-2073897,-2073894,-2073891,-2073888,-2073886,-2073883,-2073880,-2073877,-2073875,-2073872,-2073869,-2073867,-2073864,-2073861,-2073858,-2073856,-2073853,-2073850,-2073847,-2073845,-2073842,-2073839,-2073836,-2073834,-2073831,-2073828,-2073825,-2073823,-2073820,-2073817,-2073814,-2073812,-2073809,-2073806,-2073803,-2073801,-2073798,-2073795,-2073792,-2073790,-2073787,-2073784,-2073782,-2073779,-2073776,-2073773,-2073771,-2073768,-2073765,-2073762,-2073759,-2073757,-2073754,-2073751,-2073748,-2073746,-2073743,-2073740,-2073737,-2073735,-2073732,-2073729,-2073726,-2073724,-2073721,-2073718,-2073715,-2073713,-2073710,-2073707,-2073704,-2073702,-2073699,-2073696,-2073693,-2073691,-2073688,-2073685,-2073682,-2073680,-2073677,-2073674,-2073671,-2073668,-2073666,-2073663,-2073660,-2073657,-2073655,-2073652,-2073649,-2073646,-2073644,-2073641,-2073638,-2073635,-2073632,-2073630,-2073627,-2073624,-2073621,-2073619,-2073616,-2073613,-2073610,-2073608,-2073605,-2073602,-2073599,-2073596,-2073594,-2073591,-2073588,-2073585,-2073583,-2073580,-2073577,-2073574,-2073571,-2073569,-2073566,-2073563,-2073560,-2073558,-2073555,-2073552,-2073549,-2073546,-2073544,-2073541,-2073538,-2073535,-2073533,-2073530,-2073527,-2073524,-2073521,-2073519,-2073516,-2073513,-2073510,-2073507,-2073505,-2073502,-2073499,-2073496,-2073494,-2073491,-2073488,-2073485,-2073482,-2073480,-2073477,-2073474,-2073471,-2073468,-2073466,-2073463,-2073460,-2073457,-2073454,-2073452,-2073449,-2073446,-2073443,-2073440,-2073438,-2073435,-2073432,-2073429,-2073426,-2073424,-2073421,-2073418,-2073415,-2073412,-2073410,-2073407,-2073404,-2073401,-2073398,-2073396,-2073393,-2073390,-2073387,-2073384,-2073382,-2073379,-2073376,-2073373,-2073370,-2073368,-2073365,-2073362,-2073359,-2073356,-2073354,-2073351,-2073348,-2073345,-2073342,-2073340,-2073337,-2073334,-2073331,-2073328,-2073325,-2073323,-2073320,-2073317,-2073314,-2073311,-2073309,-2073306,-2073303,-2073300,-2073297,-2073294,-2073292,-2073289,-2073286,-2073283,-2073280,-2073278,-2073275,-2073272,-2073269,-2073266,-2073263,-2073261,-2073258,-2073255,-2073252,-2073249,-2073247,-2073244,-2073241,-2073238,-2073235,-2073232,-2073230,-2073227,-2073224,-2073221,-2073218,-2073215,-2073213,-2073210,-2073207,-2073204,-2073201,-2073198,-2073196,-2073193,-2073190,-2073187,-2073184,-2073182,-2073179,-2073176,-2073173,-2073170,-2073167,-2073165,-2073162,-2073159,-2073156,-2073153,-2073150,-2073148,-2073145,-2073142,-2073139,-2073136,-2073133,-2073130,-2073128,-2073125,-2073122,-2073119,-2073116,-2073113,-2073111,-2073108,-2073105,-2073102,-2073099,-2073096,-2073094,-2073091,-2073088,-2073085,-2073082,-2073079,-2073076,-2073074,-2073071,-2073068,-2073065,-2073062,-2073059,-2073057,-2073054,-2073051,-2073048,-2073045,-2073042,-2073039,-2073037,-2073034,-2073031,-2073028,-2073025,-2073022,-2073019,-2073017,-2073014,-2073011,-2073008,-2073005,-2073002,-2072999,-2072997,-2072994,-2072991,-2072988,-2072985,-2072982,-2072979,-2072977,-2072974,-2072971,-2072968,-2072965,-2072962,-2072959,-2072957,-2072954,-2072951,-2072948,-2072945,-2072942,-2072939,-2072937,-2072934,-2072931,-2072928,-2072925,-2072922,-2072919,-2072916,-2072914,-2072911,-2072908,-2072905,-2072902,-2072899,-2072896,-2072894,-2072891,-2072888,-2072885,-2072882,-2072879,-2072876,-2072873,-2072871,-2072868,-2072865,-2072862,-2072859,-2072856,-2072853,-2072850,-2072848,-2072845,-2072842,-2072839,-2072836,-2072833,-2072830,-2072827,-2072824,-2072822,-2072819,-2072816,-2072813,-2072810,-2072807,-2072804,-2072801,-2072799,-2072796,-2072793,-2072790,-2072787,-2072784,-2072781,-2072778,-2072775,-2072773,-2072770,-2072767,-2072764,-2072761,-2072758,-2072755,-2072752,-2072749,-2072747,-2072744,-2072741,-2072738,-2072735,-2072732,-2072729,-2072726,-2072723,-2072721,-2072718,-2072715,-2072712,-2072709,-2072706,-2072703,-2072700,-2072697,-2072694,-2072692,-2072689,-2072686,-2072683,-2072680,-2072677,-2072674,-2072671,-2072668,-2072665,-2072663,-2072660,-2072657,-2072654,-2072651,-2072648,-2072645,-2072642,-2072639,-2072636,-2072634,-2072631,-2072628,-2072625,-2072622,-2072619,-2072616,-2072613,-2072610,-2072607,-2072604,-2072602,-2072599,-2072596,-2072593,-2072590,-2072587,-2072584,-2072581,-2072578,-2072575,-2072572,-2072570,-2072567,-2072564,-2072561,-2072558,-2072555,-2072552,-2072549,-2072546,-2072543,-2072540,-2072537,-2072535,-2072532,-2072529,-2072526,-2072523,-2072520,-2072517,-2072514,-2072511,-2072508,-2072505,-2072502,-2072499,-2072497,-2072494,-2072491,-2072488,-2072485,-2072482,-2072479,-2072476,-2072473,-2072470,-2072467,-2072464,-2072461,-2072459,-2072456,-2072453,-2072450,-2072447,-2072444,-2072441,-2072438,-2072435,-2072432,-2072429,-2072426,-2072423,-2072420,-2072417,-2072415,-2072412,-2072409,-2072406,-2072403,-2072400,-2072397,-2072394,-2072391,-2072388,-2072385,-2072382,-2072379,-2072376,-2072373,-2072370,-2072368,-2072365,-2072362,-2072359,-2072356,-2072353,-2072350,-2072347,-2072344,-2072341,-2072338,-2072335,-2072332,-2072329,-2072326,-2072323,-2072320,-2072317,-2072315,-2072312,-2072309,-2072306,-2072303,-2072300,-2072297,-2072294,-2072291,-2072288,-2072285,-2072282,-2072279,-2072276,-2072273,-2072270,-2072267,-2072264,-2072261,-2072258,-2072256,-2072253,-2072250,-2072247,-2072244,-2072241,-2072238,-2072235,-2072232,-2072229,-2072226,-2072223,-2072220,-2072217,-2072214,-2072211,-2072208,-2072205,-2072202,-2072199,-2072196,-2072193,-2072190,-2072187,-2072184,-2072182,-2072179,-2072176,-2072173,-2072170,-2072167,-2072164,-2072161,-2072158,-2072155,-2072152,-2072149,-2072146,-2072143,-2072140,-2072137,-2072134,-2072131,-2072128,-2072125,-2072122,-2072119,-2072116,-2072113,-2072110,-2072107,-2072104,-2072101,-2072098,-2072095,-2072092,-2072089,-2072086,-2072083,-2072080,-2072077,-2072075,-2072072,-2072069,-2072066,-2072063,-2072060,-2072057,-2072054,-2072051,-2072048,-2072045,-2072042,-2072039,-2072036,-2072033,-2072030,-2072027,-2072024,-2072021,-2072018,-2072015,-2072012,-2072009,-2072006,-2072003,-2072000,-2071997,-2071994,-2071991,-2071988,-2071985,-2071982,-2071979,-2071976,-2071973,-2071970,-2071967,-2071964,-2071961,-2071958,-2071955,-2071952,-2071949,-2071946,-2071943,-2071940,-2071937,-2071934,-2071931,-2071928,-2071925,-2071922,-2071919,-2071916,-2071913,-2071910,-2071907,-2071904,-2071901,-2071898,-2071895,-2071892,-2071889,-2071886,-2071883,-2071880,-2071877,-2071874,-2071871,-2071868,-2071865,-2071862,-2071859,-2071856,-2071853,-2071850,-2071847,-2071844,-2071841,-2071838,-2071835,-2071832,-2071829,-2071826,-2071823,-2071820,-2071817,-2071814,-2071811,-2071808,-2071805,-2071802,-2071799,-2071796,-2071793,-2071790,-2071787,-2071784,-2071781,-2071778,-2071775,-2071772,-2071769,-2071766,-2071763,-2071760,-2071757,-2071754,-2071751,-2071748,-2071745,-2071741,-2071738,-2071735,-2071732,-2071729,-2071726,-2071723,-2071720,-2071717,-2071714,-2071711,-2071708,-2071705,-2071702,-2071699,-2071696,-2071693,-2071690,-2071687,-2071684,-2071681,-2071678,-2071675,-2071672,-2071669,-2071666,-2071663,-2071660,-2071657,-2071654,-2071651,-2071648,-2071645,-2071642,-2071639,-2071635,-2071632,-2071629,-2071626,-2071623,-2071620,-2071617,-2071614,-2071611,-2071608,-2071605,-2071602,-2071599,-2071596,-2071593,-2071590,-2071587,-2071584,-2071581,-2071578,-2071575,-2071572,-2071569,-2071566,-2071563,-2071559,-2071556,-2071553,-2071550,-2071547,-2071544,-2071541,-2071538,-2071535,-2071532,-2071529,-2071526,-2071523,-2071520,-2071517,-2071514,-2071511,-2071508,-2071505,-2071502,-2071499,-2071495,-2071492,-2071489,-2071486,-2071483,-2071480,-2071477,-2071474,-2071471,-2071468,-2071465,-2071462,-2071459,-2071456,-2071453,-2071450,-2071447,-2071444,-2071440,-2071437,-2071434,-2071431,-2071428,-2071425,-2071422,-2071419,-2071416,-2071413,-2071410,-2071407,-2071404,-2071401,-2071398,-2071395,-2071391,-2071388,-2071385,-2071382,-2071379,-2071376,-2071373,-2071370,-2071367,-2071364,-2071361,-2071358,-2071355,-2071352,-2071348,-2071345,-2071342,-2071339,-2071336,-2071333,-2071330,-2071327,-2071324,-2071321,-2071318,-2071315,-2071312,-2071309,-2071305,-2071302,-2071299,-2071296,-2071293,-2071290,-2071287,-2071284,-2071281,-2071278,-2071275,-2071272,-2071268,-2071265,-2071262,-2071259,-2071256,-2071253,-2071250,-2071247,-2071244,-2071241,-2071238,-2071235,-2071231,-2071228,-2071225,-2071222,-2071219,-2071216,-2071213,-2071210,-2071207,-2071204,-2071201,-2071198,-2071194,-2071191,-2071188,-2071185,-2071182,-2071179,-2071176,-2071173,-2071170,-2071167,-2071164,-2071160,-2071157,-2071154,-2071151,-2071148,-2071145,-2071142,-2071139,-2071136,-2071133,-2071129,-2071126,-2071123,-2071120,-2071117,-2071114,-2071111,-2071108,-2071105,-2071102,-2071098,-2071095,-2071092,-2071089,-2071086,-2071083,-2071080,-2071077,-2071074,-2071070,-2071067,-2071064,-2071061,-2071058,-2071055,-2071052,-2071049,-2071046,-2071043,-2071039,-2071036,-2071033,-2071030,-2071027,-2071024,-2071021,-2071018,-2071015,-2071011,-2071008,-2071005,-2071002,-2070999,-2070996,-2070993,-2070990,-2070986,-2070983,-2070980,-2070977,-2070974,-2070971,-2070968,-2070965,-2070962,-2070958,-2070955,-2070952,-2070949,-2070946,-2070943,-2070940,-2070937,-2070933,-2070930,-2070927,-2070924,-2070921,-2070918,-2070915,-2070912,-2070908,-2070905,-2070902,-2070899,-2070896,-2070893,-2070890,-2070887,-2070883,-2070880,-2070877,-2070874,-2070871,-2070868,-2070865,-2070862,-2070858,-2070855,-2070852,-2070849,-2070846,-2070843,-2070840,-2070836,-2070833,-2070830,-2070827,-2070824,-2070821,-2070818,-2070815,-2070811,-2070808,-2070805,-2070802,-2070799,-2070796,-2070793,-2070789,-2070786,-2070783,-2070780,-2070777,-2070774,-2070771,-2070767,-2070764,-2070761,-2070758,-2070755,-2070752,-2070749,-2070745,-2070742,-2070739,-2070736,-2070733,-2070730,-2070727,-2070723,-2070720,-2070717,-2070714,-2070711,-2070708,-2070704,-2070701,-2070698,-2070695,-2070692,-2070689,-2070686,-2070682,-2070679,-2070676,-2070673,-2070670,-2070667,-2070663,-2070660,-2070657,-2070654,-2070651,-2070648,-2070645,-2070641,-2070638,-2070635,-2070632,-2070629,-2070626,-2070622,-2070619,-2070616,-2070613,-2070610,-2070607,-2070603,-2070600,-2070597,-2070594,-2070591,-2070588,-2070584,-2070581,-2070578,-2070575,-2070572,-2070569,-2070565,-2070562,-2070559,-2070556,-2070553,-2070550,-2070546,-2070543,-2070540,-2070537,-2070534,-2070531,-2070527,-2070524,-2070521,-2070518,-2070515,-2070512,-2070508,-2070505,-2070502,-2070499,-2070496,-2070492,-2070489,-2070486,-2070483,-2070480,-2070477,-2070473,-2070470,-2070467,-2070464,-2070461,-2070458,-2070454,-2070451,-2070448,-2070445,-2070442,-2070438,-2070435,-2070432,-2070429,-2070426,-2070422,-2070419,-2070416,-2070413,-2070410,-2070407,-2070403,-2070400,-2070397,-2070394,-2070391,-2070387,-2070384,-2070381,-2070378,-2070375,-2070371,-2070368,-2070365,-2070362,-2070359,-2070356,-2070352,-2070349,-2070346,-2070343,-2070340,-2070336,-2070333,-2070330,-2070327,-2070324,-2070320,-2070317,-2070314,-2070311,-2070308,-2070304,-2070301,-2070298,-2070295,-2070292,-2070288,-2070285,-2070282,-2070279,-2070276,-2070272,-2070269,-2070266,-2070263,-2070260,-2070256,-2070253,-2070250,-2070247,-2070244,-2070240,-2070237,-2070234,-2070231,-2070227,-2070224,-2070221,-2070218,-2070215,-2070211,-2070208,-2070205,-2070202,-2070199,-2070195,-2070192,-2070189,-2070186,-2070183,-2070179,-2070176,-2070173,-2070170,-2070166,-2070163,-2070160,-2070157,-2070154,-2070150,-2070147,-2070144,-2070141,-2070137,-2070134,-2070131,-2070128,-2070125,-2070121,-2070118,-2070115,-2070112,-2070108,-2070105,-2070102,-2070099,-2070096,-2070092,-2070089,-2070086,-2070083,-2070079,-2070076,-2070073,-2070070,-2070067,-2070063,-2070060,-2070057,-2070054,-2070050,-2070047,-2070044,-2070041,-2070037,-2070034,-2070031,-2070028,-2070025,-2070021,-2070018,-2070015,-2070012,-2070008,-2070005,-2070002,-2069999,-2069995,-2069992,-2069989,-2069986,-2069982,-2069979,-2069976,-2069973,-2069970,-2069966,-2069963,-2069960,-2069957,-2069953,-2069950,-2069947,-2069944,-2069940,-2069937,-2069934,-2069931,-2069927,-2069924,-2069921,-2069918,-2069914,-2069911,-2069908,-2069905,-2069901,-2069898,-2069895,-2069892,-2069888,-2069885,-2069882,-2069879,-2069875,-2069872,-2069869,-2069866,-2069862,-2069859,-2069856,-2069853,-2069849,-2069846,-2069843,-2069840,-2069836,-2069833,-2069830,-2069827,-2069823,-2069820,-2069817,-2069814,-2069810,-2069807,-2069804,-2069801,-2069797,-2069794,-2069791,-2069788,-2069784,-2069781,-2069778,-2069774,-2069771,-2069768,-2069765,-2069761,-2069758,-2069755,-2069752,-2069748,-2069745,-2069742,-2069739,-2069735,-2069732,-2069729,-2069725,-2069722,-2069719,-2069716,-2069712,-2069709,-2069706,-2069703,-2069699,-2069696,-2069693,-2069690,-2069686,-2069683,-2069680,-2069676,-2069673,-2069670,-2069667,-2069663,-2069660,-2069657,-2069653,-2069650,-2069647,-2069644,-2069640,-2069637,-2069634,-2069631,-2069627,-2069624,-2069621,-2069617,-2069614,-2069611,-2069608,-2069604,-2069601,-2069598,-2069594,-2069591,-2069588,-2069585,-2069581,-2069578,-2069575,-2069571,-2069568,-2069565,-2069562,-2069558,-2069555,-2069552,-2069548,-2069545,-2069542,-2069539,-2069535,-2069532,-2069529,-2069525,-2069522,-2069519,-2069516,-2069512,-2069509,-2069506,-2069502,-2069499,-2069496,-2069492,-2069489,-2069486,-2069483,-2069479,-2069476,-2069473,-2069469,-2069466,-2069463,-2069459,-2069456,-2069453,-2069450,-2069446,-2069443,-2069440,-2069436,-2069433,-2069430,-2069426,-2069423,-2069420,-2069417,-2069413,-2069410,-2069407,-2069403,-2069400,-2069397,-2069393,-2069390,-2069387,-2069383,-2069380,-2069377,-2069374,-2069370,-2069367,-2069364,-2069360,-2069357,-2069354,-2069350,-2069347,-2069344,-2069340,-2069337,-2069334,-2069330,-2069327,-2069324,-2069321,-2069317,-2069314,-2069311,-2069307,-2069304,-2069301,-2069297,-2069294,-2069291,-2069287,-2069284,-2069281,-2069277,-2069274,-2069271,-2069267,-2069264,-2069261,-2069257,-2069254,-2069251,-2069248,-2069244,-2069241,-2069238,-2069234,-2069231,-2069228,-2069224,-2069221,-2069218,-2069214,-2069211,-2069208,-2069204,-2069201,-2069198,-2069194,-2069191,-2069188,-2069184,-2069181,-2069178,-2069174,-2069171,-2069168,-2069164,-2069161,-2069158,-2069154,-2069151,-2069148,-2069144,-2069141,-2069138,-2069134,-2069131,-2069128,-2069124,-2069121,-2069118,-2069114,-2069111,-2069108,-2069104,-2069101,-2069098,-2069094,-2069091,-2069088,-2069084,-2069081,-2069077,-2069074,-2069071,-2069067,-2069064,-2069061,-2069057,-2069054,-2069051,-2069047,-2069044,-2069041,-2069037,-2069034,-2069031,-2069027,-2069024,-2069021,-2069017,-2069014,-2069011,-2069007,-2069004,-2069000,-2068997,-2068994,-2068990,-2068987,-2068984,-2068980,-2068977,-2068974,-2068970,-2068967,-2068964,-2068960,-2068957,-2068953,-2068950,-2068947,-2068943,-2068940,-2068937,-2068933,-2068930,-2068927,-2068923,-2068920,-2068917,-2068913,-2068910,-2068906,-2068903,-2068900,-2068896,-2068893,-2068890,-2068886,-2068883,-2068880,-2068876,-2068873,-2068869,-2068866,-2068863,-2068859,-2068856,-2068853,-2068849,-2068846,-2068842,-2068839,-2068836,-2068832,-2068829,-2068826,-2068822,-2068819,-2068815,-2068812,-2068809,-2068805,-2068802,-2068799,-2068795,-2068792,-2068788,-2068785,-2068782,-2068778,-2068775,-2068772,-2068768,-2068765,-2068761,-2068758,-2068755,-2068751,-2068748,-2068745,-2068741,-2068738,-2068734,-2068731,-2068728,-2068724,-2068721,-2068717,-2068714,-2068711,-2068707,-2068704,-2068701,-2068697,-2068694,-2068690,-2068687,-2068684,-2068680,-2068677,-2068673,-2068670,-2068667,-2068663,-2068660,-2068656,-2068653,-2068650,-2068646,-2068643,-2068640,-2068636,-2068633,-2068629,-2068626,-2068623,-2068619,-2068616,-2068612,-2068609,-2068606,-2068602,-2068599,-2068595,-2068592,-2068589,-2068585,-2068582,-2068578,-2068575,-2068572,-2068568,-2068565,-2068561,-2068558,-2068555,-2068551,-2068548,-2068544,-2068541,-2068538,-2068534,-2068531,-2068527,-2068524,-2068520,-2068517,-2068514,-2068510,-2068507,-2068503,-2068500,-2068497,-2068493,-2068490,-2068486,-2068483,-2068480,-2068476,-2068473,-2068469,-2068466,-2068463,-2068459,-2068456,-2068452,-2068449,-2068445,-2068442,-2068439,-2068435,-2068432,-2068428,-2068425,-2068422,-2068418,-2068415,-2068411,-2068408,-2068404,-2068401,-2068398,-2068394,-2068391,-2068387,-2068384,-2068380,-2068377,-2068374,-2068370,-2068367,-2068363,-2068360,-2068357,-2068353,-2068350,-2068346,-2068343,-2068339,-2068336,-2068333,-2068329,-2068326,-2068322,-2068319,-2068315,-2068312,-2068309,-2068305,-2068302,-2068298,-2068295,-2068291,-2068288,-2068284,-2068281,-2068278,-2068274,-2068271,-2068267,-2068264,-2068260,-2068257,-2068254,-2068250,-2068247,-2068243,-2068240,-2068236,-2068233,-2068229,-2068226,-2068223,-2068219,-2068216,-2068212,-2068209,-2068205,-2068202,-2068199,-2068195,-2068192,-2068188,-2068185,-2068181,-2068178,-2068174,-2068171,-2068168,-2068164,-2068161,-2068157,-2068154,-2068150,-2068147,-2068143,-2068140,-2068136,-2068133,-2068130,-2068126,-2068123,-2068119,-2068116,-2068112,-2068109,-2068105,-2068102,-2068098,-2068095,-2068092,-2068088,-2068085,-2068081,-2068078,-2068074,-2068071,-2068067,-2068064,-2068060,-2068057,-2068054,-2068050,-2068047,-2068043,-2068040,-2068036,-2068033,-2068029,-2068026,-2068022,-2068019,-2068015,-2068012,-2068009,-2068005,-2068002,-2067998,-2067995,-2067991,-2067988,-2067984,-2067981,-2067977,-2067974,-2067970,-2067967,-2067963,-2067960,-2067957,-2067953,-2067950,-2067946,-2067943,-2067939,-2067936,-2067932,-2067929,-2067925,-2067922,-2067918,-2067915,-2067911,-2067908,-2067904,-2067901,-2067897,-2067894,-2067891,-2067887,-2067884,-2067880,-2067877,-2067873,-2067870,-2067866,-2067863,-2067859,-2067856,-2067852,-2067849,-2067845,-2067842,-2067838,-2067835,-2067831,-2067828,-2067824,-2067821,-2067817,-2067814,-2067810,-2067807,-2067803,-2067800,-2067796,-2067793,-2067790,-2067786,-2067783,-2067779,-2067776,-2067772,-2067769,-2067765,-2067762,-2067758,-2067755,-2067751,-2067748,-2067744,-2067741,-2067737,-2067734,-2067730,-2067727,-2067723,-2067720,-2067716,-2067713,-2067709,-2067706,-2067702,-2067699,-2067695,-2067692,-2067688,-2067685,-2067681,-2067678,-2067674,-2067671,-2067667,-2067664,-2067660,-2067657,-2067653,-2067650,-2067646,-2067643,-2067639,-2067636,-2067632,-2067629,-2067625,-2067622,-2067618,-2067615,-2067611,-2067608,-2067604,-2067601,-2067597,-2067594,-2067590,-2067587,-2067583,-2067579,-2067576,-2067572,-2067569,-2067565,-2067562,-2067558,-2067555,-2067551,-2067548,-2067544,-2067541,-2067537,-2067534,-2067530,-2067527,-2067523,-2067520,-2067516,-2067513,-2067509,-2067506,-2067502,-2067499,-2067495,-2067492,-2067488,-2067485,-2067481,-2067477,-2067474,-2067470,-2067467,-2067463,-2067460,-2067456,-2067453,-2067449,-2067446,-2067442,-2067439,-2067435,-2067432,-2067428,-2067425,-2067421,-2067418,-2067414,-2067410,-2067407,-2067403,-2067400,-2067396,-2067393,-2067389,-2067386,-2067382,-2067379,-2067375,-2067372,-2067368,-2067365,-2067361,-2067357,-2067354,-2067350,-2067347,-2067343,-2067340,-2067336,-2067333,-2067329,-2067326,-2067322,-2067319,-2067315,-2067311,-2067308,-2067304,-2067301,-2067297,-2067294,-2067290,-2067287,-2067283,-2067280,-2067276,-2067272,-2067269,-2067265,-2067262,-2067258,-2067255,-2067251,-2067248,-2067244,-2067241,-2067237,-2067233,-2067230,-2067226,-2067223,-2067219,-2067216,-2067212,-2067209,-2067205,-2067202,-2067198,-2067194,-2067191,-2067187,-2067184,-2067180,-2067177,-2067173,-2067170,-2067166,-2067162,-2067159,-2067155,-2067152,-2067148,-2067145,-2067141,-2067137,-2067134,-2067130,-2067127,-2067123,-2067120,-2067116,-2067113,-2067109,-2067105,-2067102,-2067098,-2067095,-2067091,-2067088,-2067084,-2067080,-2067077,-2067073,-2067070,-2067066,-2067063,-2067059,-2067056,-2067052,-2067048,-2067045,-2067041,-2067038,-2067034,-2067031,-2067027,-2067023,-2067020,-2067016,-2067013,-2067009,-2067006,-2067002,-2066998,-2066995,-2066991,-2066988,-2066984,-2066980,-2066977,-2066973,-2066970,-2066966,-2066963,-2066959,-2066955,-2066952,-2066948,-2066945,-2066941,-2066938,-2066934,-2066930,-2066927,-2066923,-2066920,-2066916,-2066912,-2066909,-2066905,-2066902,-2066898,-2066895,-2066891,-2066887,-2066884,-2066880,-2066877,-2066873,-2066869,-2066866,-2066862,-2066859,-2066855,-2066851,-2066848,-2066844,-2066841,-2066837,-2066833,-2066830,-2066826,-2066823,-2066819,-2066816,-2066812,-2066808,-2066805,-2066801,-2066798,-2066794,-2066790,-2066787,-2066783,-2066780,-2066776,-2066772,-2066769,-2066765,-2066762,-2066758,-2066754,-2066751,-2066747,-2066744,-2066740,-2066736,-2066733,-2066729,-2066726,-2066722,-2066718,-2066715,-2066711,-2066708,-2066704,-2066700,-2066697,-2066693,-2066689,-2066686,-2066682,-2066679,-2066675,-2066671,-2066668,-2066664,-2066661,-2066657,-2066653,-2066650,-2066646,-2066643,-2066639,-2066635,-2066632,-2066628,-2066624,-2066621,-2066617,-2066614,-2066610,-2066606,-2066603,-2066599,-2066596,-2066592,-2066588,-2066585,-2066581,-2066577,-2066574,-2066570,-2066567,-2066563,-2066559,-2066556,-2066552,-2066548,-2066545,-2066541,-2066538,-2066534,-2066530,-2066527,-2066523,-2066519,-2066516,-2066512,-2066509,-2066505,-2066501,-2066498,-2066494,-2066490,-2066487,-2066483,-2066480,-2066476,-2066472,-2066469,-2066465,-2066461,-2066458,-2066454,-2066451,-2066447,-2066443,-2066440,-2066436,-2066432,-2066429,-2066425,-2066421,-2066418,-2066414,-2066411,-2066407,-2066403,-2066400,-2066396,-2066392,-2066389,-2066385,-2066381,-2066378,-2066374,-2066370,-2066367,-2066363,-2066360,-2066356,-2066352,-2066349,-2066345,-2066341,-2066338,-2066334,-2066330,-2066327,-2066323,-2066319,-2066316,-2066312,-2066309,-2066305,-2066301,-2066298,-2066294,-2066290,-2066287,-2066283,-2066279,-2066276,-2066272,-2066268,-2066265,-2066261,-2066257,-2066254,-2066250,-2066246,-2066243,-2066239,-2066235,-2066232,-2066228,-2066225,-2066221,-2066217,-2066214,-2066210,-2066206,-2066203,-2066199,-2066195,-2066192,-2066188,-2066184,-2066181,-2066177,-2066173,-2066170,-2066166,-2066162,-2066159,-2066155,-2066151,-2066148,-2066144,-2066140,-2066137,-2066133,-2066129,-2066126,-2066122,-2066118,-2066115,-2066111,-2066107,-2066104,-2066100,-2066096,-2066093,-2066089,-2066085,-2066082,-2066078,-2066074,-2066071,-2066067,-2066063,-2066060,-2066056,-2066052,-2066049,-2066045,-2066041,-2066037,-2066034,-2066030,-2066026,-2066023,-2066019,-2066015,-2066012,-2066008,-2066004,-2066001,-2065997,-2065993,-2065990,-2065986,-2065982,-2065979,-2065975,-2065971,-2065968,-2065964,-2065960,-2065957,-2065953,-2065949,-2065945,-2065942,-2065938,-2065934,-2065931,-2065927,-2065923,-2065920,-2065916,-2065912,-2065909,-2065905,-2065901,-2065898,-2065894,-2065890,-2065886,-2065883,-2065879,-2065875,-2065872,-2065868,-2065864,-2065861,-2065857,-2065853,-2065849,-2065846,-2065842,-2065838,-2065835,-2065831,-2065827,-2065824,-2065820,-2065816,-2065813,-2065809,-2065805,-2065801,-2065798,-2065794,-2065790,-2065787,-2065783,-2065779,-2065775,-2065772,-2065768,-2065764,-2065761,-2065757,-2065753,-2065750,-2065746,-2065742,-2065738,-2065735,-2065731,-2065727,-2065724,-2065720,-2065716,-2065712,-2065709,-2065705,-2065701,-2065698,-2065694,-2065690,-2065686,-2065683,-2065679,-2065675,-2065672,-2065668,-2065664,-2065660,-2065657,-2065653,-2065649,-2065646,-2065642,-2065638,-2065634,-2065631,-2065627,-2065623,-2065620,-2065616,-2065612,-2065608,-2065605,-2065601,-2065597,-2065594,-2065590,-2065586,-2065582,-2065579,-2065575,-2065571,-2065567,-2065564,-2065560,-2065556,-2065553,-2065549,-2065545,-2065541,-2065538,-2065534,-2065530,-2065526,-2065523,-2065519,-2065515,-2065512,-2065508,-2065504,-2065500,-2065497,-2065493,-2065489,-2065485,-2065482,-2065478,-2065474,-2065470,-2065467,-2065463,-2065459,-2065456,-2065452,-2065448,-2065444,-2065441,-2065437,-2065433,-2065429,-2065426,-2065422,-2065418,-2065414,-2065411,-2065407,-2065403,-2065399,-2065396,-2065392,-2065388,-2065384,-2065381,-2065377,-2065373,-2065369,-2065366,-2065362,-2065358,-2065354,-2065351,-2065347,-2065343,-2065339,-2065336,-2065332,-2065328,-2065324,-2065321,-2065317,-2065313,-2065309,-2065306,-2065302,-2065298,-2065294,-2065291,-2065287,-2065283,-2065279,-2065276,-2065272,-2065268,-2065264,-2065261,-2065257,-2065253,-2065249,-2065246,-2065242,-2065238,-2065234,-2065231,-2065227,-2065223,-2065219,-2065216,-2065212,-2065208,-2065204,-2065201,-2065197,-2065193,-2065189,-2065185,-2065182,-2065178,-2065174,-2065170,-2065167,-2065163,-2065159,-2065155,-2065152,-2065148,-2065144,-2065140,-2065136,-2065133,-2065129,-2065125,-2065121,-2065118,-2065114,-2065110,-2065106,-2065103,-2065099,-2065095,-2065091,-2065087,-2065084,-2065080,-2065076,-2065072,-2065069,-2065065,-2065061,-2065057,-2065053,-2065050,-2065046,-2065042,-2065038,-2065035,-2065031,-2065027,-2065023,-2065019,-2065016,-2065012,-2065008,-2065004,-2065001,-2064997,-2064993,-2064989,-2064985,-2064982,-2064978,-2064974,-2064970,-2064966,-2064963,-2064959,-2064955,-2064951,-2064948,-2064944,-2064940,-2064936,-2064932,-2064929,-2064925,-2064921,-2064917,-2064913,-2064910,-2064906,-2064902,-2064898,-2064894,-2064891,-2064887,-2064883,-2064879,-2064875,-2064872,-2064868,-2064864,-2064860,-2064856,-2064853,-2064849,-2064845,-2064841,-2064837,-2064834,-2064830,-2064826,-2064822,-2064818,-2064815,-2064811,-2064807,-2064803,-2064799,-2064796,-2064792,-2064788,-2064784,-2064780,-2064777,-2064773,-2064769,-2064765,-2064761,-2064758,-2064754,-2064750,-2064746,-2064742,-2064739,-2064735,-2064731,-2064727,-2064723,-2064719,-2064716,-2064712,-2064708,-2064704,-2064700,-2064697,-2064693,-2064689,-2064685,-2064681,-2064678,-2064674,-2064670,-2064666,-2064662,-2064658,-2064655,-2064651,-2064647,-2064643,-2064639,-2064636,-2064632,-2064628,-2064624,-2064620,-2064616,-2064613,-2064609,-2064605,-2064601,-2064597,-2064593,-2064590,-2064586,-2064582,-2064578,-2064574,-2064571,-2064567,-2064563,-2064559,-2064555,-2064551,-2064548,-2064544,-2064540,-2064536,-2064532,-2064528,-2064525,-2064521,-2064517,-2064513,-2064509,-2064505,-2064502,-2064498,-2064494,-2064490,-2064486,-2064482,-2064479,-2064475,-2064471,-2064467,-2064463,-2064459,-2064456,-2064452,-2064448,-2064444,-2064440,-2064436,-2064433,-2064429,-2064425,-2064421,-2064417,-2064413,-2064409,-2064406,-2064402,-2064398,-2064394,-2064390,-2064386,-2064383,-2064379,-2064375,-2064371,-2064367,-2064363,-2064359,-2064356,-2064352,-2064348,-2064344,-2064340,-2064336,-2064333,-2064329,-2064325,-2064321,-2064317,-2064313,-2064309,-2064306,-2064302,-2064298,-2064294,-2064290,-2064286,-2064282,-2064279,-2064275,-2064271,-2064267,-2064263,-2064259,-2064255,-2064252,-2064248,-2064244,-2064240,-2064236,-2064232,-2064228,-2064225,-2064221,-2064217,-2064213,-2064209,-2064205,-2064201,-2064198,-2064194,-2064190,-2064186,-2064182,-2064178,-2064174,-2064170,-2064167,-2064163,-2064159,-2064155,-2064151,-2064147,-2064143,-2064140,-2064136,-2064132,-2064128,-2064124,-2064120,-2064116,-2064112,-2064109,-2064105,-2064101,-2064097,-2064093,-2064089,-2064085,-2064081,-2064078,-2064074,-2064070,-2064066,-2064062,-2064058,-2064054,-2064050,-2064047,-2064043,-2064039,-2064035,-2064031,-2064027,-2064023,-2064019,-2064015,-2064012,-2064008,-2064004,-2064000,-2063996,-2063992,-2063988,-2063984,-2063981,-2063977,-2063973,-2063969,-2063965,-2063961,-2063957,-2063953,-2063949,-2063946,-2063942,-2063938,-2063934,-2063930,-2063926,-2063922,-2063918,-2063914,-2063911,-2063907,-2063903,-2063899,-2063895,-2063891,-2063887,-2063883,-2063879,-2063875,-2063872,-2063868,-2063864,-2063860,-2063856,-2063852,-2063848,-2063844,-2063840,-2063836,-2063833,-2063829,-2063825,-2063821,-2063817,-2063813,-2063809,-2063805,-2063801,-2063797,-2063794,-2063790,-2063786,-2063782,-2063778,-2063774,-2063770,-2063766,-2063762,-2063758,-2063755,-2063751,-2063747,-2063743,-2063739,-2063735,-2063731,-2063727,-2063723,-2063719,-2063715,-2063711,-2063708,-2063704,-2063700,-2063696,-2063692,-2063688,-2063684,-2063680,-2063676,-2063672,-2063668,-2063665,-2063661,-2063657,-2063653,-2063649,-2063645,-2063641,-2063637,-2063633,-2063629,-2063625,-2063621,-2063617,-2063614,-2063610,-2063606,-2063602,-2063598,-2063594,-2063590,-2063586,-2063582,-2063578,-2063574,-2063570,-2063566,-2063563,-2063559,-2063555,-2063551,-2063547,-2063543,-2063539,-2063535,-2063531,-2063527,-2063523,-2063519,-2063515,-2063511,-2063508,-2063504,-2063500,-2063496,-2063492,-2063488,-2063484,-2063480,-2063476,-2063472,-2063468,-2063464,-2063460,-2063456,-2063452,-2063449,-2063445,-2063441,-2063437,-2063433,-2063429,-2063425,-2063421,-2063417,-2063413,-2063409,-2063405,-2063401,-2063397,-2063393,-2063389,-2063385,-2063382,-2063378,-2063374,-2063370,-2063366,-2063362,-2063358,-2063354,-2063350,-2063346,-2063342,-2063338,-2063334,-2063330,-2063326,-2063322,-2063318,-2063314,-2063310,-2063307,-2063303,-2063299,-2063295,-2063291,-2063287,-2063283,-2063279,-2063275,-2063271,-2063267,-2063263,-2063259,-2063255,-2063251,-2063247,-2063243,-2063239,-2063235,-2063231,-2063227,-2063223,-2063219,-2063216,-2063212,-2063208,-2063204,-2063200,-2063196,-2063192,-2063188,-2063184,-2063180,-2063176,-2063172,-2063168,-2063164,-2063160,-2063156,-2063152,-2063148,-2063144,-2063140,-2063136,-2063132,-2063128,-2063124,-2063120,-2063116,-2063112,-2063108,-2063104,-2063101,-2063097,-2063093,-2063089,-2063085,-2063081,-2063077,-2063073,-2063069,-2063065,-2063061,-2063057,-2063053,-2063049,-2063045,-2063041,-2063037,-2063033,-2063029,-2063025,-2063021,-2063017,-2063013,-2063009,-2063005,-2063001,-2062997,-2062993,-2062989,-2062985,-2062981,-2062977,-2062973,-2062969,-2062965,-2062961,-2062957,-2062953,-2062949,-2062945,-2062941,-2062937,-2062933,-2062929,-2062925,-2062921,-2062917,-2062913,-2062909,-2062905,-2062901,-2062897,-2062893,-2062889,-2062885,-2062881,-2062877,-2062874,-2062870,-2062866,-2062862,-2062858,-2062854,-2062850,-2062846,-2062842,-2062838,-2062834,-2062830,-2062826,-2062822,-2062818,-2062814,-2062810,-2062806,-2062802,-2062798,-2062794,-2062790,-2062786,-2062782,-2062778,-2062774,-2062770,-2062766,-2062762,-2062758,-2062754,-2062750,-2062746,-2062742,-2062738,-2062734,-2062729,-2062725,-2062721,-2062717,-2062713,-2062709,-2062705,-2062701,-2062697,-2062693,-2062689,-2062685,-2062681,-2062677,-2062673,-2062669,-2062665,-2062661,-2062657,-2062653,-2062649,-2062645,-2062641,-2062637,-2062633,-2062629,-2062625,-2062621,-2062617,-2062613,-2062609,-2062605,-2062601,-2062597,-2062593,-2062589,-2062585,-2062581,-2062577,-2062573,-2062569,-2062565,-2062561,-2062557,-2062553,-2062549,-2062545,-2062541,-2062537,-2062533,-2062529,-2062525,-2062521,-2062517,-2062513,-2062509,-2062504,-2062500,-2062496,-2062492,-2062488,-2062484,-2062480,-2062476,-2062472,-2062468,-2062464,-2062460,-2062456,-2062452,-2062448,-2062444,-2062440,-2062436,-2062432,-2062428,-2062424,-2062420,-2062416,-2062412,-2062408,-2062404,-2062400,-2062396,-2062392,-2062387,-2062383,-2062379,-2062375,-2062371,-2062367,-2062363,-2062359,-2062355,-2062351,-2062347,-2062343,-2062339,-2062335,-2062331,-2062327,-2062323,-2062319,-2062315,-2062311,-2062307,-2062303,-2062299,-2062294,-2062290,-2062286,-2062282,-2062278,-2062274,-2062270,-2062266,-2062262,-2062258,-2062254,-2062250,-2062246,-2062242,-2062238,-2062234,-2062230,-2062226,-2062222,-2062217,-2062213,-2062209,-2062205,-2062201,-2062197,-2062193,-2062189,-2062185,-2062181,-2062177,-2062173,-2062169,-2062165,-2062161,-2062157,-2062153,-2062148,-2062144,-2062140,-2062136,-2062132,-2062128,-2062124,-2062120,-2062116,-2062112,-2062108,-2062104,-2062100,-2062096,-2062092,-2062087,-2062083,-2062079,-2062075,-2062071,-2062067,-2062063,-2062059,-2062055,-2062051,-2062047,-2062043,-2062039,-2062035,-2062031,-2062026,-2062022,-2062018,-2062014,-2062010,-2062006,-2062002,-2061998,-2061994,-2061990,-2061986,-2061982,-2061978,-2061973,-2061969,-2061965,-2061961,-2061957,-2061953,-2061949,-2061945,-2061941,-2061937,-2061933,-2061929,-2061924,-2061920,-2061916,-2061912,-2061908,-2061904,-2061900,-2061896,-2061892,-2061888,-2061884,-2061880,-2061875,-2061871,-2061867,-2061863,-2061859,-2061855,-2061851,-2061847,-2061843,-2061839,-2061835,-2061830,-2061826,-2061822,-2061818,-2061814,-2061810,-2061806,-2061802,-2061798,-2061794,-2061789,-2061785,-2061781,-2061777,-2061773,-2061769,-2061765,-2061761,-2061757,-2061753,-2061749,-2061744,-2061740,-2061736,-2061732,-2061728,-2061724,-2061720,-2061716,-2061712,-2061707,-2061703,-2061699,-2061695,-2061691,-2061687,-2061683,-2061679,-2061675,-2061671,-2061666,-2061662,-2061658,-2061654,-2061650,-2061646,-2061642,-2061638,-2061634,-2061629,-2061625,-2061621,-2061617,-2061613,-2061609,-2061605,-2061601,-2061597,-2061592,-2061588,-2061584,-2061580,-2061576,-2061572,-2061568,-2061564,-2061560,-2061555,-2061551,-2061547,-2061543,-2061539,-2061535,-2061531,-2061527,-2061522,-2061518,-2061514,-2061510,-2061506,-2061502,-2061498,-2061494,-2061489,-2061485,-2061481,-2061477,-2061473,-2061469,-2061465,-2061461,-2061456,-2061452,-2061448,-2061444,-2061440,-2061436,-2061432,-2061428,-2061423,-2061419,-2061415,-2061411,-2061407,-2061403,-2061399,-2061394,-2061390,-2061386,-2061382,-2061378,-2061374,-2061370,-2061366,-2061361,-2061357,-2061353,-2061349,-2061345,-2061341,-2061337,-2061332,-2061328,-2061324,-2061320,-2061316,-2061312,-2061308,-2061303,-2061299,-2061295,-2061291,-2061287,-2061283,-2061279,-2061274,-2061270,-2061266,-2061262,-2061258,-2061254,-2061250,-2061245,-2061241,-2061237,-2061233,-2061229,-2061225,-2061221,-2061216,-2061212,-2061208,-2061204,-2061200,-2061196,-2061192,-2061187,-2061183,-2061179,-2061175,-2061171,-2061167,-2061162,-2061158,-2061154,-2061150,-2061146,-2061142,-2061138,-2061133,-2061129,-2061125,-2061121,-2061117,-2061113,-2061108,-2061104,-2061100,-2061096,-2061092,-2061088,-2061083,-2061079,-2061075,-2061071,-2061067,-2061063,-2061058,-2061054,-2061050,-2061046,-2061042,-2061038,-2061033,-2061029,-2061025,-2061021,-2061017,-2061013,-2061008,-2061004,-2061000,-2060996,-2060992,-2060988,-2060983,-2060979,-2060975,-2060971,-2060967,-2060963,-2060958,-2060954,-2060950,-2060946,-2060942,-2060938,-2060933,-2060929,-2060925,-2060921,-2060917,-2060912,-2060908,-2060904,-2060900,-2060896,-2060892,-2060887,-2060883,-2060879,-2060875,-2060871,-2060867,-2060862,-2060858,-2060854,-2060850,-2060846,-2060841,-2060837,-2060833,-2060829,-2060825,-2060820,-2060816,-2060812,-2060808,-2060804,-2060800,-2060795,-2060791,-2060787,-2060783,-2060779,-2060774,-2060770,-2060766,-2060762,-2060758,-2060753,-2060749,-2060745,-2060741,-2060737,-2060733,-2060728,-2060724,-2060720,-2060716,-2060712,-2060707,-2060703,-2060699,-2060695,-2060691,-2060686,-2060682,-2060678,-2060674,-2060670,-2060665,-2060661,-2060657,-2060653,-2060649,-2060644,-2060640,-2060636,-2060632,-2060628,-2060623,-2060619,-2060615,-2060611,-2060607,-2060602,-2060598,-2060594,-2060590,-2060585,-2060581,-2060577,-2060573,-2060569,-2060564,-2060560,-2060556,-2060552,-2060548,-2060543,-2060539,-2060535,-2060531,-2060527,-2060522,-2060518,-2060514,-2060510,-2060505,-2060501,-2060497,-2060493,-2060489,-2060484,-2060480,-2060476,-2060472,-2060468,-2060463,-2060459,-2060455,-2060451,-2060446,-2060442,-2060438,-2060434,-2060430,-2060425,-2060421,-2060417,-2060413,-2060408,-2060404,-2060400,-2060396,-2060392,-2060387,-2060383,-2060379,-2060375,-2060370,-2060366,-2060362,-2060358,-2060353,-2060349,-2060345,-2060341,-2060337,-2060332,-2060328,-2060324,-2060320,-2060315,-2060311,-2060307,-2060303,-2060298,-2060294,-2060290,-2060286,-2060282,-2060277,-2060273,-2060269,-2060265,-2060260,-2060256,-2060252,-2060248,-2060243,-2060239,-2060235,-2060231,-2060226,-2060222,-2060218,-2060214,-2060210,-2060205,-2060201,-2060197,-2060193,-2060188,-2060184,-2060180,-2060176,-2060171,-2060167,-2060163,-2060159,-2060154,-2060150,-2060146,-2060142,-2060137,-2060133,-2060129,-2060125,-2060120,-2060116,-2060112,-2060108,-2060103,-2060099,-2060095,-2060091,-2060086,-2060082,-2060078,-2060074,-2060069,-2060065,-2060061,-2060057,-2060052,-2060048,-2060044,-2060040,-2060035,-2060031,-2060027,-2060023,-2060018,-2060014,-2060010,-2060005,-2060001,-2059997,-2059993,-2059988,-2059984,-2059980,-2059976,-2059971,-2059967,-2059963,-2059959,-2059954,-2059950,-2059946,-2059942,-2059937,-2059933,-2059929,-2059924,-2059920,-2059916,-2059912,-2059907,-2059903,-2059899,-2059895,-2059890,-2059886,-2059882,-2059878,-2059873,-2059869,-2059865,-2059860,-2059856,-2059852,-2059848,-2059843,-2059839,-2059835,-2059831,-2059826,-2059822,-2059818,-2059813,-2059809,-2059805,-2059801,-2059796,-2059792,-2059788,-2059783,-2059779,-2059775,-2059771,-2059766,-2059762,-2059758,-2059753,-2059749,-2059745,-2059741,-2059736,-2059732,-2059728,-2059723,-2059719,-2059715,-2059711,-2059706,-2059702,-2059698,-2059693,-2059689,-2059685,-2059681,-2059676,-2059672,-2059668,-2059663,-2059659,-2059655,-2059651,-2059646,-2059642,-2059638,-2059633,-2059629,-2059625,-2059621,-2059616,-2059612,-2059608,-2059603,-2059599,-2059595,-2059590,-2059586,-2059582,-2059578,-2059573,-2059569,-2059565,-2059560,-2059556,-2059552,-2059547,-2059543,-2059539,-2059535,-2059530,-2059526,-2059522,-2059517,-2059513,-2059509,-2059504,-2059500,-2059496,-2059492,-2059487,-2059483,-2059479,-2059474,-2059470,-2059466,-2059461,-2059457,-2059453,-2059448,-2059444,-2059440,-2059436,-2059431,-2059427,-2059423,-2059418,-2059414,-2059410,-2059405,-2059401,-2059397,-2059392,-2059388,-2059384,-2059379,-2059375,-2059371,-2059367,-2059362,-2059358,-2059354,-2059349,-2059345,-2059341,-2059336,-2059332,-2059328,-2059323,-2059319,-2059315,-2059310,-2059306,-2059302,-2059297,-2059293,-2059289,-2059284,-2059280,-2059276,-2059271,-2059267,-2059263,-2059258,-2059254,-2059250,-2059245,-2059241,-2059237,-2059233,-2059228,-2059224,-2059220,-2059215,-2059211,-2059207,-2059202,-2059198,-2059194,-2059189,-2059185,-2059181,-2059176,-2059172,-2059168,-2059163,-2059159,-2059155,-2059150,-2059146,-2059142,-2059137,-2059133,-2059129,-2059124,-2059120,-2059115,-2059111,-2059107,-2059102,-2059098,-2059094,-2059089,-2059085,-2059081,-2059076,-2059072,-2059068,-2059063,-2059059,-2059055,-2059050,-2059046,-2059042,-2059037,-2059033,-2059029,-2059024,-2059020,-2059016,-2059011,-2059007,-2059003,-2058998,-2058994,-2058990,-2058985,-2058981,-2058976,-2058972,-2058968,-2058963,-2058959,-2058955,-2058950,-2058946,-2058942,-2058937,-2058933,-2058929,-2058924,-2058920,-2058915,-2058911,-2058907,-2058902,-2058898,-2058894,-2058889,-2058885,-2058881,-2058876,-2058872,-2058868,-2058863,-2058859,-2058854,-2058850,-2058846,-2058841,-2058837,-2058833,-2058828,-2058824,-2058820,-2058815,-2058811,-2058806,-2058802,-2058798,-2058793,-2058789,-2058785,-2058780,-2058776,-2058772,-2058767,-2058763,-2058758,-2058754,-2058750,-2058745,-2058741,-2058737,-2058732,-2058728,-2058723,-2058719,-2058715,-2058710,-2058706,-2058702,-2058697,-2058693,-2058688,-2058684,-2058680,-2058675,-2058671,-2058667,-2058662,-2058658,-2058653,-2058649,-2058645,-2058640,-2058636,-2058632,-2058627,-2058623,-2058618,-2058614,-2058610,-2058605,-2058601,-2058596,-2058592,-2058588,-2058583,-2058579,-2058575,-2058570,-2058566,-2058561,-2058557,-2058553,-2058548,-2058544,-2058539,-2058535,-2058531,-2058526,-2058522,-2058517,-2058513,-2058509,-2058504,-2058500,-2058495,-2058491,-2058487,-2058482,-2058478,-2058474,-2058469,-2058465,-2058460,-2058456,-2058452,-2058447,-2058443,-2058438,-2058434,-2058430,-2058425,-2058421,-2058416,-2058412,-2058408,-2058403,-2058399,-2058394,-2058390,-2058386,-2058381,-2058377,-2058372,-2058368,-2058364,-2058359,-2058355,-2058350,-2058346,-2058341,-2058337,-2058333,-2058328,-2058324,-2058319,-2058315,-2058311,-2058306,-2058302,-2058297,-2058293,-2058289,-2058284,-2058280,-2058275,-2058271,-2058267,-2058262,-2058258,-2058253,-2058249,-2058244,-2058240,-2058236,-2058231,-2058227,-2058222,-2058218,-2058214,-2058209,-2058205,-2058200,-2058196,-2058191,-2058187,-2058183,-2058178,-2058174,-2058169,-2058165,-2058160,-2058156,-2058152,-2058147,-2058143,-2058138,-2058134,-2058130,-2058125,-2058121,-2058116,-2058112,-2058107,-2058103,-2058099,-2058094,-2058090,-2058085,-2058081,-2058076,-2058072,-2058068,-2058063,-2058059,-2058054,-2058050,-2058045,-2058041,-2058037,-2058032,-2058028,-2058023,-2058019,-2058014,-2058010,-2058005,-2058001,-2057997,-2057992,-2057988,-2057983,-2057979,-2057974,-2057970,-2057966,-2057961,-2057957,-2057952,-2057948,-2057943,-2057939,-2057934,-2057930,-2057926,-2057921,-2057917,-2057912,-2057908,-2057903,-2057899,-2057894,-2057890,-2057886,-2057881,-2057877,-2057872,-2057868,-2057863,-2057859,-2057854,-2057850,-2057846,-2057841,-2057837,-2057832,-2057828,-2057823,-2057819,-2057814,-2057810,-2057805,-2057801,-2057797,-2057792,-2057788,-2057783,-2057779,-2057774,-2057770,-2057765,-2057761,-2057756,-2057752,-2057748,-2057743,-2057739,-2057734,-2057730,-2057725,-2057721,-2057716,-2057712,-2057707,-2057703,-2057698,-2057694,-2057690,-2057685,-2057681,-2057676,-2057672,-2057667,-2057663,-2057658,-2057654,-2057649,-2057645,-2057640,-2057636,-2057631,-2057627,-2057623,-2057618,-2057614,-2057609,-2057605,-2057600,-2057596,-2057591,-2057587,-2057582,-2057578,-2057573,-2057569,-2057564,-2057560,-2057555,-2057551,-2057547,-2057542,-2057538,-2057533,-2057529,-2057524,-2057520,-2057515,-2057511,-2057506,-2057502,-2057497,-2057493,-2057488,-2057484,-2057479,-2057475,-2057470,-2057466,-2057461,-2057457,-2057452,-2057448,-2057443,-2057439,-2057435,-2057430,-2057426,-2057421,-2057417,-2057412,-2057408,-2057403,-2057399,-2057394,-2057390,-2057385,-2057381,-2057376,-2057372,-2057367,-2057363,-2057358,-2057354,-2057349,-2057345,-2057340,-2057336,-2057331,-2057327,-2057322,-2057318,-2057313,-2057309,-2057304,-2057300,-2057295,-2057291,-2057286,-2057282,-2057277,-2057273,-2057268,-2057264,-2057259,-2057255,-2057250,-2057246,-2057241,-2057237,-2057232,-2057228,-2057223,-2057219,-2057214,-2057210,-2057205,-2057201,-2057196,-2057192,-2057187,-2057183,-2057178,-2057174,-2057169,-2057165,-2057160,-2057156,-2057151,-2057147,-2057142,-2057138,-2057133,-2057129,-2057124,-2057120,-2057115,-2057111,-2057106,-2057102,-2057097,-2057093,-2057088,-2057084,-2057079,-2057075,-2057070,-2057065,-2057061,-2057056,-2057052,-2057047,-2057043,-2057038,-2057034,-2057029,-2057025,-2057020,-2057016,-2057011,-2057007,-2057002,-2056998,-2056993,-2056989,-2056984,-2056980,-2056975,-2056971,-2056966,-2056962,-2056957,-2056952,-2056948,-2056943,-2056939,-2056934,-2056930,-2056925,-2056921,-2056916,-2056912,-2056907,-2056903,-2056898,-2056894,-2056889,-2056885,-2056880,-2056875,-2056871,-2056866,-2056862,-2056857,-2056853,-2056848,-2056844,-2056839,-2056835,-2056830,-2056826,-2056821,-2056817,-2056812,-2056807,-2056803,-2056798,-2056794,-2056789,-2056785,-2056780,-2056776,-2056771,-2056767,-2056762,-2056757,-2056753,-2056748,-2056744,-2056739,-2056735,-2056730,-2056726,-2056721,-2056717,-2056712,-2056708,-2056703,-2056698,-2056694,-2056689,-2056685,-2056680,-2056676,-2056671,-2056667,-2056662,-2056657,-2056653,-2056648,-2056644,-2056639,-2056635,-2056630,-2056626,-2056621,-2056617,-2056612,-2056607,-2056603,-2056598,-2056594,-2056589,-2056585,-2056580,-2056575,-2056571,-2056566,-2056562,-2056557,-2056553,-2056548,-2056544,-2056539,-2056534,-2056530,-2056525,-2056521,-2056516,-2056512,-2056507,-2056503,-2056498,-2056493,-2056489,-2056484,-2056480,-2056475,-2056471,-2056466,-2056461,-2056457,-2056452,-2056448,-2056443,-2056439,-2056434,-2056429,-2056425,-2056420,-2056416,-2056411,-2056407,-2056402,-2056397,-2056393,-2056388,-2056384,-2056379,-2056375,-2056370,-2056365,-2056361,-2056356,-2056352,-2056347,-2056343,-2056338,-2056333,-2056329,-2056324,-2056320,-2056315,-2056311,-2056306,-2056301,-2056297,-2056292,-2056288,-2056283,-2056278,-2056274,-2056269,-2056265,-2056260,-2056256,-2056251,-2056246,-2056242,-2056237,-2056233,-2056228,-2056223,-2056219,-2056214,-2056210,-2056205,-2056200,-2056196,-2056191,-2056187,-2056182,-2056178,-2056173,-2056168,-2056164,-2056159,-2056155,-2056150,-2056145,-2056141,-2056136,-2056132,-2056127,-2056122,-2056118,-2056113,-2056109,-2056104,-2056099,-2056095,-2056090,-2056086,-2056081,-2056076,-2056072,-2056067,-2056063,-2056058,-2056053,-2056049,-2056044,-2056040,-2056035,-2056030,-2056026,-2056021,-2056017,-2056012,-2056007,-2056003,-2055998,-2055994,-2055989,-2055984,-2055980,-2055975,-2055971,-2055966,-2055961,-2055957,-2055952,-2055948,-2055943,-2055938,-2055934,-2055929,-2055924,-2055920,-2055915,-2055911,-2055906,-2055901,-2055897,-2055892,-2055888,-2055883,-2055878,-2055874,-2055869,-2055864,-2055860,-2055855,-2055851,-2055846,-2055841,-2055837,-2055832,-2055828,-2055823,-2055818,-2055814,-2055809,-2055804,-2055800,-2055795,-2055791,-2055786,-2055781,-2055777,-2055772,-2055767,-2055763,-2055758,-2055754,-2055749,-2055744,-2055740,-2055735,-2055730,-2055726,-2055721,-2055717,-2055712,-2055707,-2055703,-2055698,-2055693,-2055689,-2055684,-2055680,-2055675,-2055670,-2055666,-2055661,-2055656,-2055652,-2055647,-2055642,-2055638,-2055633,-2055629,-2055624,-2055619,-2055615,-2055610,-2055605,-2055601,-2055596,-2055591,-2055587,-2055582,-2055578,-2055573,-2055568,-2055564,-2055559,-2055554,-2055550,-2055545,-2055540,-2055536,-2055531,-2055526,-2055522,-2055517,-2055513,-2055508,-2055503,-2055499,-2055494,-2055489,-2055485,-2055480,-2055475,-2055471,-2055466,-2055461,-2055457,-2055452,-2055447,-2055443,-2055438,-2055433,-2055429,-2055424,-2055420,-2055415,-2055410,-2055406,-2055401,-2055396,-2055392,-2055387,-2055382,-2055378,-2055373,-2055368,-2055364,-2055359,-2055354,-2055350,-2055345,-2055340,-2055336,-2055331,-2055326,-2055322,-2055317,-2055312,-2055308,-2055303,-2055298,-2055294,-2055289,-2055284,-2055280,-2055275,-2055270,-2055266,-2055261,-2055256,-2055252,-2055247,-2055242,-2055238,-2055233,-2055228,-2055224,-2055219,-2055214,-2055210,-2055205,-2055200,-2055196,-2055191,-2055186,-2055182,-2055177,-2055172,-2055168,-2055163,-2055158,-2055154,-2055149,-2055144,-2055140,-2055135,-2055130,-2055126,-2055121,-2055116,-2055112,-2055107,-2055102,-2055098,-2055093,-2055088,-2055083,-2055079,-2055074,-2055069,-2055065,-2055060,-2055055,-2055051,-2055046,-2055041,-2055037,-2055032,-2055027,-2055023,-2055018,-2055013,-2055009,-2055004,-2054999,-2054994,-2054990,-2054985,-2054980,-2054976,-2054971,-2054966,-2054962,-2054957,-2054952,-2054948,-2054943,-2054938,-2054933,-2054929,-2054924,-2054919,-2054915,-2054910,-2054905,-2054901,-2054896,-2054891,-2054887,-2054882,-2054877,-2054872,-2054868,-2054863,-2054858,-2054854,-2054849,-2054844,-2054840,-2054835,-2054830,-2054825,-2054821,-2054816,-2054811,-2054807,-2054802,-2054797,-2054793,-2054788,-2054783,-2054778,-2054774,-2054769,-2054764,-2054760,-2054755,-2054750,-2054745,-2054741,-2054736,-2054731,-2054727,-2054722,-2054717,-2054712,-2054708,-2054703,-2054698,-2054694,-2054689,-2054684,-2054679,-2054675,-2054670,-2054665,-2054661,-2054656,-2054651,-2054646,-2054642,-2054637,-2054632,-2054628,-2054623,-2054618,-2054613,-2054609,-2054604,-2054599,-2054595,-2054590,-2054585,-2054580,-2054576,-2054571,-2054566,-2054562,-2054557,-2054552,-2054547,-2054543,-2054538,-2054533,-2054528,-2054524,-2054519,-2054514,-2054510,-2054505,-2054500,-2054495,-2054491,-2054486,-2054481,-2054476,-2054472,-2054467,-2054462,-2054458,-2054453,-2054448,-2054443,-2054439,-2054434,-2054429,-2054424,-2054420,-2054415,-2054410,-2054405,-2054401,-2054396,-2054391,-2054386,-2054382,-2054377,-2054372,-2054368,-2054363,-2054358,-2054353,-2054349,-2054344,-2054339,-2054334,-2054330,-2054325,-2054320,-2054315,-2054311,-2054306,-2054301,-2054296,-2054292,-2054287,-2054282,-2054277,-2054273,-2054268,-2054263,-2054258,-2054254,-2054249,-2054244,-2054239,-2054235,-2054230,-2054225,-2054220,-2054216,-2054211,-2054206,-2054201,-2054197,-2054192,-2054187,-2054182,-2054178,-2054173,-2054168,-2054163,-2054159,-2054154,-2054149,-2054144,-2054140,-2054135,-2054130,-2054125,-2054121,-2054116,-2054111,-2054106,-2054102,-2054097,-2054092,-2054087,-2054083,-2054078,-2054073,-2054068,-2054063,-2054059,-2054054,-2054049,-2054044,-2054040,-2054035,-2054030,-2054025,-2054021,-2054016,-2054011,-2054006,-2054002,-2053997,-2053992,-2053987,-2053982,-2053978,-2053973,-2053968,-2053963,-2053959,-2053954,-2053949,-2053944,-2053939,-2053935,-2053930,-2053925,-2053920,-2053916,-2053911,-2053906,-2053901,-2053897,-2053892,-2053887,-2053882,-2053877,-2053873,-2053868,-2053863,-2053858,-2053853,-2053849,-2053844,-2053839,-2053834,-2053830,-2053825,-2053820,-2053815,-2053810,-2053806,-2053801,-2053796,-2053791,-2053787,-2053782,-2053777,-2053772,-2053767,-2053763,-2053758,-2053753,-2053748,-2053743,-2053739,-2053734,-2053729,-2053724,-2053720,-2053715,-2053710,-2053705,-2053700,-2053696,-2053691,-2053686,-2053681,-2053676,-2053672,-2053667,-2053662,-2053657,-2053652,-2053648,-2053643,-2053638,-2053633,-2053628,-2053624,-2053619,-2053614,-2053609,-2053604,-2053600,-2053595,-2053590,-2053585,-2053580,-2053576,-2053571,-2053566,-2053561,-2053556,-2053552,-2053547,-2053542,-2053537,-2053532,-2053528,-2053523,-2053518,-2053513,-2053508,-2053504,-2053499,-2053494,-2053489,-2053484,-2053479,-2053475,-2053470,-2053465,-2053460,-2053455,-2053451,-2053446,-2053441,-2053436,-2053431,-2053427,-2053422,-2053417,-2053412,-2053407,-2053402,-2053398,-2053393,-2053388,-2053383,-2053378,-2053374,-2053369,-2053364,-2053359,-2053354,-2053349,-2053345,-2053340,-2053335,-2053330,-2053325,-2053321,-2053316,-2053311,-2053306,-2053301,-2053296,-2053292,-2053287,-2053282,-2053277,-2053272,-2053267,-2053263,-2053258,-2053253,-2053248,-2053243,-2053238,-2053234,-2053229,-2053224,-2053219,-2053214,-2053210,-2053205,-2053200,-2053195,-2053190,-2053185,-2053181,-2053176,-2053171,-2053166,-2053161,-2053156,-2053152,-2053147,-2053142,-2053137,-2053132,-2053127,-2053122,-2053118,-2053113,-2053108,-2053103,-2053098,-2053093,-2053089,-2053084,-2053079,-2053074,-2053069,-2053064,-2053060,-2053055,-2053050,-2053045,-2053040,-2053035,-2053030,-2053026,-2053021,-2053016,-2053011,-2053006,-2053001,-2052997,-2052992,-2052987,-2052982,-2052977,-2052972,-2052967,-2052963,-2052958,-2052953,-2052948,-2052943,-2052938,-2052933,-2052929,-2052924,-2052919,-2052914,-2052909,-2052904,-2052900,-2052895,-2052890,-2052885,-2052880,-2052875,-2052870,-2052866,-2052861,-2052856,-2052851,-2052846,-2052841,-2052836,-2052831,-2052827,-2052822,-2052817,-2052812,-2052807,-2052802,-2052797,-2052793,-2052788,-2052783,-2052778,-2052773,-2052768,-2052763,-2052759,-2052754,-2052749,-2052744,-2052739,-2052734,-2052729,-2052724,-2052720,-2052715,-2052710,-2052705,-2052700,-2052695,-2052690,-2052685,-2052681,-2052676,-2052671,-2052666,-2052661,-2052656,-2052651,-2052646,-2052642,-2052637,-2052632,-2052627,-2052622,-2052617,-2052612,-2052607,-2052603,-2052598,-2052593,-2052588,-2052583,-2052578,-2052573,-2052568,-2052564,-2052559,-2052554,-2052549,-2052544,-2052539,-2052534,-2052529,-2052524,-2052520,-2052515,-2052510,-2052505,-2052500,-2052495,-2052490,-2052485,-2052480,-2052476,-2052471,-2052466,-2052461,-2052456,-2052451,-2052446,-2052441,-2052436,-2052432,-2052427,-2052422,-2052417,-2052412,-2052407,-2052402,-2052397,-2052392,-2052388,-2052383,-2052378,-2052373,-2052368,-2052363,-2052358,-2052353,-2052348,-2052343,-2052339,-2052334,-2052329,-2052324,-2052319,-2052314,-2052309,-2052304,-2052299,-2052294,-2052290,-2052285,-2052280,-2052275,-2052270,-2052265,-2052260,-2052255,-2052250,-2052245,-2052240,-2052236,-2052231,-2052226,-2052221,-2052216,-2052211,-2052206,-2052201,-2052196,-2052191,-2052186,-2052182,-2052177,-2052172,-2052167,-2052162,-2052157,-2052152,-2052147,-2052142,-2052137,-2052132,-2052128,-2052123,-2052118,-2052113,-2052108,-2052103,-2052098,-2052093,-2052088,-2052083,-2052078,-2052073,-2052068,-2052064,-2052059,-2052054,-2052049,-2052044,-2052039,-2052034,-2052029,-2052024,-2052019,-2052014,-2052009,-2052004,-2052000,-2051995,-2051990,-2051985,-2051980,-2051975,-2051970,-2051965,-2051960,-2051955,-2051950,-2051945,-2051940,-2051935,-2051931,-2051926,-2051921,-2051916,-2051911,-2051906,-2051901,-2051896,-2051891,-2051886,-2051881,-2051876,-2051871,-2051866,-2051861,-2051857,-2051852,-2051847,-2051842,-2051837,-2051832,-2051827,-2051822,-2051817,-2051812,-2051807,-2051802,-2051797,-2051792,-2051787,-2051782,-2051778,-2051773,-2051768,-2051763,-2051758,-2051753,-2051748,-2051743,-2051738,-2051733,-2051728,-2051723,-2051718,-2051713,-2051708,-2051703,-2051698,-2051693,-2051688,-2051684,-2051679,-2051674,-2051669,-2051664,-2051659,-2051654,-2051649,-2051644,-2051639,-2051634,-2051629,-2051624,-2051619,-2051614,-2051609,-2051604,-2051599,-2051594,-2051589,-2051584,-2051579,-2051575,-2051570,-2051565,-2051560,-2051555,-2051550,-2051545,-2051540,-2051535,-2051530,-2051525,-2051520,-2051515,-2051510,-2051505,-2051500,-2051495,-2051490,-2051485,-2051480,-2051475,-2051470,-2051465,-2051460,-2051455,-2051450,-2051445,-2051440,-2051436,-2051431,-2051426,-2051421,-2051416,-2051411,-2051406,-2051401,-2051396,-2051391,-2051386,-2051381,-2051376,-2051371,-2051366,-2051361,-2051356,-2051351,-2051346,-2051341,-2051336,-2051331,-2051326,-2051321,-2051316,-2051311,-2051306,-2051301,-2051296,-2051291,-2051286,-2051281,-2051276,-2051271,-2051266,-2051261,-2051256,-2051251,-2051246,-2051241,-2051236,-2051231,-2051226,-2051221,-2051216,-2051211,-2051207,-2051202,-2051197,-2051192,-2051187,-2051182,-2051177,-2051172,-2051167,-2051162,-2051157,-2051152,-2051147,-2051142,-2051137,-2051132,-2051127,-2051122,-2051117,-2051112,-2051107,-2051102,-2051097,-2051092,-2051087,-2051082,-2051077,-2051072,-2051067,-2051062,-2051057,-2051052,-2051047,-2051042,-2051037,-2051032,-2051027,-2051022,-2051017,-2051012,-2051007,-2051002,-2050997,-2050992,-2050987,-2050982,-2050977,-2050972,-2050967,-2050962,-2050957,-2050952,-2050947,-2050942,-2050937,-2050932,-2050927,-2050922,-2050917,-2050912,-2050907,-2050902,-2050897,-2050892,-2050887,-2050882,-2050877,-2050872,-2050866,-2050861,-2050856,-2050851,-2050846,-2050841,-2050836,-2050831,-2050826,-2050821,-2050816,-2050811,-2050806,-2050801,-2050796,-2050791,-2050786,-2050781,-2050776,-2050771,-2050766,-2050761,-2050756,-2050751,-2050746,-2050741,-2050736,-2050731,-2050726,-2050721,-2050716,-2050711,-2050706,-2050701,-2050696,-2050691,-2050686,-2050681,-2050676,-2050671,-2050666,-2050661,-2050656,-2050651,-2050646,-2050641,-2050635,-2050630,-2050625,-2050620,-2050615,-2050610,-2050605,-2050600,-2050595,-2050590,-2050585,-2050580,-2050575,-2050570,-2050565,-2050560,-2050555,-2050550,-2050545,-2050540,-2050535,-2050530,-2050525,-2050520,-2050515,-2050510,-2050505,-2050500,-2050494,-2050489,-2050484,-2050479,-2050474,-2050469,-2050464,-2050459,-2050454,-2050449,-2050444,-2050439,-2050434,-2050429,-2050424,-2050419,-2050414,-2050409,-2050404,-2050399,-2050394,-2050389,-2050383,-2050378,-2050373,-2050368,-2050363,-2050358,-2050353,-2050348,-2050343,-2050338,-2050333,-2050328,-2050323,-2050318,-2050313,-2050308,-2050303,-2050298,-2050293,-2050287,-2050282,-2050277,-2050272,-2050267,-2050262,-2050257,-2050252,-2050247,-2050242,-2050237,-2050232,-2050227,-2050222,-2050217,-2050212,-2050207,-2050201,-2050196,-2050191,-2050186,-2050181,-2050176,-2050171,-2050166,-2050161,-2050156,-2050151,-2050146,-2050141,-2050136,-2050131,-2050125,-2050120,-2050115,-2050110,-2050105,-2050100,-2050095,-2050090,-2050085,-2050080,-2050075,-2050070,-2050065,-2050060,-2050054,-2050049,-2050044,-2050039,-2050034,-2050029,-2050024,-2050019,-2050014,-2050009,-2050004,-2049999,-2049994,-2049988,-2049983,-2049978,-2049973,-2049968,-2049963,-2049958,-2049953,-2049948,-2049943,-2049938,-2049933,-2049927,-2049922,-2049917,-2049912,-2049907,-2049902,-2049897,-2049892,-2049887,-2049882,-2049877,-2049872,-2049866,-2049861,-2049856,-2049851,-2049846,-2049841,-2049836,-2049831,-2049826,-2049821,-2049816,-2049810,-2049805,-2049800,-2049795,-2049790,-2049785,-2049780,-2049775,-2049770,-2049765,-2049759,-2049754,-2049749,-2049744,-2049739,-2049734,-2049729,-2049724,-2049719,-2049714,-2049709,-2049703,-2049698,-2049693,-2049688,-2049683,-2049678,-2049673,-2049668,-2049663,-2049657,-2049652,-2049647,-2049642,-2049637,-2049632,-2049627,-2049622,-2049617,-2049612,-2049606,-2049601,-2049596,-2049591,-2049586,-2049581,-2049576,-2049571,-2049566,-2049560,-2049555,-2049550,-2049545,-2049540,-2049535,-2049530,-2049525,-2049520,-2049514,-2049509,-2049504,-2049499,-2049494,-2049489,-2049484,-2049479,-2049473,-2049468,-2049463,-2049458,-2049453,-2049448,-2049443,-2049438,-2049433,-2049427,-2049422,-2049417,-2049412,-2049407,-2049402,-2049397,-2049392,-2049386,-2049381,-2049376,-2049371,-2049366,-2049361,-2049356,-2049351,-2049345,-2049340,-2049335,-2049330,-2049325,-2049320,-2049315,-2049310,-2049304,-2049299,-2049294,-2049289,-2049284,-2049279,-2049274,-2049268,-2049263,-2049258,-2049253,-2049248,-2049243,-2049238,-2049233,-2049227,-2049222,-2049217,-2049212,-2049207,-2049202,-2049197,-2049191,-2049186,-2049181,-2049176,-2049171,-2049166,-2049161,-2049155,-2049150,-2049145,-2049140,-2049135,-2049130,-2049125,-2049119,-2049114,-2049109,-2049104,-2049099,-2049094,-2049089,-2049083,-2049078,-2049073,-2049068,-2049063,-2049058,-2049053,-2049047,-2049042,-2049037,-2049032,-2049027,-2049022,-2049016,-2049011,-2049006,-2049001,-2048996,-2048991,-2048986,-2048980,-2048975,-2048970,-2048965,-2048960,-2048955,-2048949,-2048944,-2048939,-2048934,-2048929,-2048924,-2048919,-2048913,-2048908,-2048903,-2048898,-2048893,-2048888,-2048882,-2048877,-2048872,-2048867,-2048862,-2048857,-2048851,-2048846,-2048841,-2048836,-2048831,-2048826,-2048820,-2048815,-2048810,-2048805,-2048800,-2048795,-2048789,-2048784,-2048779,-2048774,-2048769,-2048764,-2048758,-2048753,-2048748,-2048743,-2048738,-2048733,-2048727,-2048722,-2048717,-2048712,-2048707,-2048702,-2048696,-2048691,-2048686,-2048681,-2048676,-2048670,-2048665,-2048660,-2048655,-2048650,-2048645,-2048639,-2048634,-2048629,-2048624,-2048619,-2048613,-2048608,-2048603,-2048598,-2048593,-2048588,-2048582,-2048577,-2048572,-2048567,-2048562,-2048556,-2048551,-2048546,-2048541,-2048536,-2048531,-2048525,-2048520,-2048515,-2048510,-2048505,-2048499,-2048494,-2048489,-2048484,-2048479,-2048473,-2048468,-2048463,-2048458,-2048453,-2048447,-2048442,-2048437,-2048432,-2048427,-2048422,-2048416,-2048411,-2048406,-2048401,-2048396,-2048390,-2048385,-2048380,-2048375,-2048370,-2048364,-2048359,-2048354,-2048349,-2048344,-2048338,-2048333,-2048328,-2048323,-2048318,-2048312,-2048307,-2048302,-2048297,-2048291,-2048286,-2048281,-2048276,-2048271,-2048265,-2048260,-2048255,-2048250,-2048245,-2048239,-2048234,-2048229,-2048224,-2048219,-2048213,-2048208,-2048203,-2048198,-2048193,-2048187,-2048182,-2048177,-2048172,-2048166,-2048161,-2048156,-2048151,-2048146,-2048140,-2048135,-2048130,-2048125,-2048120,-2048114,-2048109,-2048104,-2048099,-2048093,-2048088,-2048083,-2048078,-2048073,-2048067,-2048062,-2048057,-2048052,-2048046,-2048041,-2048036,-2048031,-2048026,-2048020,-2048015,-2048010,-2048005,-2047999,-2047994,-2047989,-2047984,-2047978,-2047973,-2047968,-2047963,-2047958,-2047952,-2047947,-2047942,-2047937,-2047931,-2047926,-2047921,-2047916,-2047911,-2047905,-2047900,-2047895,-2047890,-2047884,-2047879,-2047874,-2047869,-2047863,-2047858,-2047853,-2047848,-2047842,-2047837,-2047832,-2047827,-2047821,-2047816,-2047811,-2047806,-2047801,-2047795,-2047790,-2047785,-2047780,-2047774,-2047769,-2047764,-2047759,-2047753,-2047748,-2047743,-2047738,-2047732,-2047727,-2047722,-2047717,-2047711,-2047706,-2047701,-2047696,-2047690,-2047685,-2047680,-2047675,-2047669,-2047664,-2047659,-2047654,-2047648,-2047643,-2047638,-2047633,-2047627,-2047622,-2047617,-2047612,-2047606,-2047601,-2047596,-2047591,-2047585,-2047580,-2047575,-2047570,-2047564,-2047559,-2047554,-2047549,-2047543,-2047538,-2047533,-2047527,-2047522,-2047517,-2047512,-2047506,-2047501,-2047496,-2047491,-2047485,-2047480,-2047475,-2047470,-2047464,-2047459,-2047454,-2047449,-2047443,-2047438,-2047433,-2047427,-2047422,-2047417,-2047412,-2047406,-2047401,-2047396,-2047391,-2047385,-2047380,-2047375,-2047369,-2047364,-2047359,-2047354,-2047348,-2047343,-2047338,-2047333,-2047327,-2047322,-2047317,-2047311,-2047306,-2047301,-2047296,-2047290,-2047285,-2047280,-2047275,-2047269,-2047264,-2047259,-2047253,-2047248,-2047243,-2047238,-2047232,-2047227,-2047222,-2047216,-2047211,-2047206,-2047201,-2047195,-2047190,-2047185,-2047179,-2047174,-2047169,-2047164,-2047158,-2047153,-2047148,-2047142,-2047137,-2047132,-2047127,-2047121,-2047116,-2047111,-2047105,-2047100,-2047095,-2047090,-2047084,-2047079,-2047074,-2047068,-2047063,-2047058,-2047052,-2047047,-2047042,-2047037,-2047031,-2047026,-2047021,-2047015,-2047010,-2047005,-2047000,-2046994,-2046989,-2046984,-2046978,-2046973,-2046968,-2046962,-2046957,-2046952,-2046947,-2046941,-2046936,-2046931,-2046925,-2046920,-2046915,-2046909,-2046904,-2046899,-2046893,-2046888,-2046883,-2046878,-2046872,-2046867,-2046862,-2046856,-2046851,-2046846,-2046840,-2046835,-2046830,-2046824,-2046819,-2046814,-2046809,-2046803,-2046798,-2046793,-2046787,-2046782,-2046777,-2046771,-2046766,-2046761,-2046755,-2046750,-2046745,-2046739,-2046734,-2046729,-2046723,-2046718,-2046713,-2046707,-2046702,-2046697,-2046692,-2046686,-2046681,-2046676,-2046670,-2046665,-2046660,-2046654,-2046649,-2046644,-2046638,-2046633,-2046628,-2046622,-2046617,-2046612,-2046606,-2046601,-2046596,-2046590,-2046585,-2046580,-2046574,-2046569,-2046564,-2046558,-2046553,-2046548,-2046542,-2046537,-2046532,-2046526,-2046521,-2046516,-2046510,-2046505,-2046500,-2046494,-2046489,-2046484,-2046478,-2046473,-2046468,-2046462,-2046457,-2046452,-2046446,-2046441,-2046436,-2046430,-2046425,-2046420,-2046414,-2046409,-2046404,-2046398,-2046393,-2046388,-2046382,-2046377,-2046372,-2046366,-2046361,-2046356,-2046350,-2046345,-2046340,-2046334,-2046329,-2046323,-2046318,-2046313,-2046307,-2046302,-2046297,-2046291,-2046286,-2046281,-2046275,-2046270,-2046265,-2046259,-2046254,-2046249,-2046243,-2046238,-2046233,-2046227,-2046222,-2046216,-2046211,-2046206,-2046200,-2046195,-2046190,-2046184,-2046179,-2046174,-2046168,-2046163,-2046158,-2046152,-2046147,-2046141,-2046136,-2046131,-2046125,-2046120,-2046115,-2046109,-2046104,-2046099,-2046093,-2046088,-2046082,-2046077,-2046072,-2046066,-2046061,-2046056,-2046050,-2046045,-2046040,-2046034,-2046029,-2046023,-2046018,-2046013,-2046007,-2046002,-2045997,-2045991,-2045986,-2045980,-2045975,-2045970,-2045964,-2045959,-2045954,-2045948,-2045943,-2045938,-2045932,-2045927,-2045921,-2045916,-2045911,-2045905,-2045900,-2045895,-2045889,-2045884,-2045878,-2045873,-2045868,-2045862,-2045857,-2045851,-2045846,-2045841,-2045835,-2045830,-2045825,-2045819,-2045814,-2045808,-2045803,-2045798,-2045792,-2045787,-2045781,-2045776,-2045771,-2045765,-2045760,-2045755,-2045749,-2045744,-2045738,-2045733,-2045728,-2045722,-2045717,-2045711,-2045706,-2045701,-2045695,-2045690,-2045684,-2045679,-2045674,-2045668,-2045663,-2045658,-2045652,-2045647,-2045641,-2045636,-2045631,-2045625,-2045620,-2045614,-2045609,-2045604,-2045598,-2045593,-2045587,-2045582,-2045577,-2045571,-2045566,-2045560,-2045555,-2045550,-2045544,-2045539,-2045533,-2045528,-2045523,-2045517,-2045512,-2045506,-2045501,-2045496,-2045490,-2045485,-2045479,-2045474,-2045468,-2045463,-2045458,-2045452,-2045447,-2045441,-2045436,-2045431,-2045425,-2045420,-2045414,-2045409,-2045404,-2045398,-2045393,-2045387,-2045382,-2045377,-2045371,-2045366,-2045360,-2045355,-2045349,-2045344,-2045339,-2045333,-2045328,-2045322,-2045317,-2045312,-2045306,-2045301,-2045295,-2045290,-2045284,-2045279,-2045274,-2045268,-2045263,-2045257,-2045252,-2045246,-2045241,-2045236,-2045230,-2045225,-2045219,-2045214,-2045208,-2045203,-2045198,-2045192,-2045187,-2045181,-2045176,-2045170,-2045165,-2045160,-2045154,-2045149,-2045143,-2045138,-2045132,-2045127,-2045122,-2045116,-2045111,-2045105,-2045100,-2045094,-2045089,-2045084,-2045078,-2045073,-2045067,-2045062,-2045056,-2045051,-2045046,-2045040,-2045035,-2045029,-2045024,-2045018,-2045013,-2045007,-2045002,-2044997,-2044991,-2044986,-2044980,-2044975,-2044969,-2044964,-2044958,-2044953,-2044948,-2044942,-2044937,-2044931,-2044926,-2044920,-2044915,-2044909,-2044904,-2044899,-2044893,-2044888,-2044882,-2044877,-2044871,-2044866,-2044860,-2044855,-2044850,-2044844,-2044839,-2044833,-2044828,-2044822,-2044817,-2044811,-2044806,-2044800,-2044795,-2044790,-2044784,-2044779,-2044773,-2044768,-2044762,-2044757,-2044751,-2044746,-2044740,-2044735,-2044730,-2044724,-2044719,-2044713,-2044708,-2044702,-2044697,-2044691,-2044686,-2044680,-2044675,-2044669,-2044664,-2044659,-2044653,-2044648,-2044642,-2044637,-2044631,-2044626,-2044620,-2044615,-2044609,-2044604,-2044598,-2044593,-2044587,-2044582,-2044577,-2044571,-2044566,-2044560,-2044555,-2044549,-2044544,-2044538,-2044533,-2044527,-2044522,-2044516,-2044511,-2044505,-2044500,-2044494,-2044489,-2044483,-2044478,-2044473,-2044467,-2044462,-2044456,-2044451,-2044445,-2044440,-2044434,-2044429,-2044423,-2044418,-2044412,-2044407,-2044401,-2044396,-2044390,-2044385,-2044379,-2044374,-2044368,-2044363,-2044357,-2044352,-2044346,-2044341,-2044335,-2044330,-2044325,-2044319,-2044314,-2044308,-2044303,-2044297,-2044292,-2044286,-2044281,-2044275,-2044270,-2044264,-2044259,-2044253,-2044248,-2044242,-2044237,-2044231,-2044226,-2044220,-2044215,-2044209,-2044204,-2044198,-2044193,-2044187,-2044182,-2044176,-2044171,-2044165,-2044160,-2044154,-2044149,-2044143,-2044138,-2044132,-2044127,-2044121,-2044116,-2044110,-2044105,-2044099,-2044094,-2044088,-2044083,-2044077,-2044072,-2044066,-2044061,-2044055,-2044050,-2044044,-2044039,-2044033,-2044028,-2044022,-2044017,-2044011,-2044006,-2044000,-2043995,-2043989,-2043984,-2043978,-2043973,-2043967,-2043962,-2043956,-2043950,-2043945,-2043939,-2043934,-2043928,-2043923,-2043917,-2043912,-2043906,-2043901,-2043895,-2043890,-2043884,-2043879,-2043873,-2043868,-2043862,-2043857,-2043851,-2043846,-2043840,-2043835,-2043829,-2043824,-2043818,-2043813,-2043807,-2043801,-2043796,-2043790,-2043785,-2043779,-2043774,-2043768,-2043763,-2043757,-2043752,-2043746,-2043741,-2043735,-2043730,-2043724,-2043719,-2043713,-2043708,-2043702,-2043696,-2043691,-2043685,-2043680,-2043674,-2043669,-2043663,-2043658,-2043652,-2043647,-2043641,-2043636,-2043630,-2043625,-2043619,-2043613,-2043608,-2043602,-2043597,-2043591,-2043586,-2043580,-2043575,-2043569,-2043564,-2043558,-2043553,-2043547,-2043541,-2043536,-2043530,-2043525,-2043519,-2043514,-2043508,-2043503,-2043497,-2043492,-2043486,-2043480,-2043475,-2043469,-2043464,-2043458,-2043453,-2043447,-2043442,-2043436,-2043431,-2043425,-2043419,-2043414,-2043408,-2043403,-2043397,-2043392,-2043386,-2043381,-2043375,-2043369,-2043364,-2043358,-2043353,-2043347,-2043342,-2043336,-2043331,-2043325,-2043320,-2043314,-2043308,-2043303,-2043297,-2043292,-2043286,-2043281,-2043275,-2043269,-2043264,-2043258,-2043253,-2043247,-2043242,-2043236,-2043231,-2043225,-2043219,-2043214,-2043208,-2043203,-2043197,-2043192,-2043186,-2043180,-2043175,-2043169,-2043164,-2043158,-2043153,-2043147,-2043141,-2043136,-2043130,-2043125,-2043119,-2043114,-2043108,-2043103,-2043097,-2043091,-2043086,-2043080,-2043075,-2043069,-2043063,-2043058,-2043052,-2043047,-2043041,-2043036,-2043030,-2043024,-2043019,-2043013,-2043008,-2043002,-2042997,-2042991,-2042985,-2042980,-2042974,-2042969,-2042963,-2042958,-2042952,-2042946,-2042941,-2042935,-2042930,-2042924,-2042918,-2042913,-2042907,-2042902,-2042896,-2042891,-2042885,-2042879,-2042874,-2042868,-2042863,-2042857,-2042851,-2042846,-2042840,-2042835,-2042829,-2042823,-2042818,-2042812,-2042807,-2042801,-2042796,-2042790,-2042784,-2042779,-2042773,-2042768,-2042762,-2042756,-2042751,-2042745,-2042740,-2042734,-2042728,-2042723,-2042717,-2042712,-2042706,-2042700,-2042695,-2042689,-2042684,-2042678,-2042672,-2042667,-2042661,-2042656,-2042650,-2042644,-2042639,-2042633,-2042628,-2042622,-2042616,-2042611,-2042605,-2042600,-2042594,-2042588,-2042583,-2042577,-2042572,-2042566,-2042560,-2042555,-2042549,-2042543,-2042538,-2042532,-2042527,-2042521,-2042515,-2042510,-2042504,-2042499,-2042493,-2042487,-2042482,-2042476,-2042471,-2042465,-2042459,-2042454,-2042448,-2042442,-2042437,-2042431,-2042426,-2042420,-2042414,-2042409,-2042403,-2042397,-2042392,-2042386,-2042381,-2042375,-2042369,-2042364,-2042358,-2042353,-2042347,-2042341,-2042336,-2042330,-2042324,-2042319,-2042313,-2042308,-2042302,-2042296,-2042291,-2042285,-2042279,-2042274,-2042268,-2042263,-2042257,-2042251,-2042246,-2042240,-2042234,-2042229,-2042223,-2042217,-2042212,-2042206,-2042201,-2042195,-2042189,-2042184,-2042178,-2042172,-2042167,-2042161,-2042156,-2042150,-2042144,-2042139,-2042133,-2042127,-2042122,-2042116,-2042110,-2042105,-2042099,-2042093,-2042088,-2042082,-2042077,-2042071,-2042065,-2042060,-2042054,-2042048,-2042043,-2042037,-2042031,-2042026,-2042020,-2042015,-2042009,-2042003,-2041998,-2041992,-2041986,-2041981,-2041975,-2041969,-2041964,-2041958,-2041952,-2041947,-2041941,-2041935,-2041930,-2041924,-2041918,-2041913,-2041907,-2041902,-2041896,-2041890,-2041885,-2041879,-2041873,-2041868,-2041862,-2041856,-2041851,-2041845,-2041839,-2041834,-2041828,-2041822,-2041817,-2041811,-2041805,-2041800,-2041794,-2041788,-2041783,-2041777,-2041771,-2041766,-2041760,-2041754,-2041749,-2041743,-2041737,-2041732,-2041726,-2041720,-2041715,-2041709,-2041703,-2041698,-2041692,-2041686,-2041681,-2041675,-2041669,-2041664,-2041658,-2041652,-2041647,-2041641,-2041635,-2041630,-2041624,-2041618,-2041613,-2041607,-2041601,-2041596,-2041590,-2041584,-2041579,-2041573,-2041567,-2041562,-2041556,-2041550,-2041545,-2041539,-2041533,-2041528,-2041522,-2041516,-2041511,-2041505,-2041499,-2041494,-2041488,-2041482,-2041477,-2041471,-2041465,-2041459,-2041454,-2041448,-2041442,-2041437,-2041431,-2041425,-2041420,-2041414,-2041408,-2041403,-2041397,-2041391,-2041386,-2041380,-2041374,-2041368,-2041363,-2041357,-2041351,-2041346,-2041340,-2041334,-2041329,-2041323,-2041317,-2041312,-2041306,-2041300,-2041295,-2041289,-2041283,-2041277,-2041272,-2041266,-2041260,-2041255,-2041249,-2041243,-2041238,-2041232,-2041226,-2041220,-2041215,-2041209,-2041203,-2041198,-2041192,-2041186,-2041181,-2041175,-2041169,-2041163,-2041158,-2041152,-2041146,-2041141,-2041135,-2041129,-2041124,-2041118,-2041112,-2041106,-2041101,-2041095,-2041089,-2041084,-2041078,-2041072,-2041066,-2041061,-2041055,-2041049,-2041044,-2041038,-2041032,-2041027,-2041021,-2041015,-2041009,-2041004,-2040998,-2040992,-2040987,-2040981,-2040975,-2040969,-2040964,-2040958,-2040952,-2040947,-2040941,-2040935,-2040929,-2040924,-2040918,-2040912,-2040906,-2040901,-2040895,-2040889,-2040884,-2040878,-2040872,-2040866,-2040861,-2040855,-2040849,-2040844,-2040838,-2040832,-2040826,-2040821,-2040815,-2040809,-2040803,-2040798,-2040792,-2040786,-2040781,-2040775,-2040769,-2040763,-2040758,-2040752,-2040746,-2040740,-2040735,-2040729,-2040723,-2040718,-2040712,-2040706,-2040700,-2040695,-2040689,-2040683,-2040677,-2040672,-2040666,-2040660,-2040654,-2040649,-2040643,-2040637,-2040632,-2040626,-2040620,-2040614,-2040609,-2040603,-2040597,-2040591,-2040586,-2040580,-2040574,-2040568,-2040563,-2040557,-2040551,-2040545,-2040540,-2040534,-2040528,-2040522,-2040517,-2040511,-2040505,-2040499,-2040494,-2040488,-2040482,-2040476,-2040471,-2040465,-2040459,-2040454,-2040448,-2040442,-2040436,-2040431,-2040425,-2040419,-2040413,-2040407,-2040402,-2040396,-2040390,-2040384,-2040379,-2040373,-2040367,-2040361,-2040356,-2040350,-2040344,-2040338,-2040333,-2040327,-2040321,-2040315,-2040310,-2040304,-2040298,-2040292,-2040287,-2040281,-2040275,-2040269,-2040264,-2040258,-2040252,-2040246,-2040241,-2040235,-2040229,-2040223,-2040217,-2040212,-2040206,-2040200,-2040194,-2040189,-2040183,-2040177,-2040171,-2040166,-2040160,-2040154,-2040148,-2040143,-2040137,-2040131,-2040125,-2040119,-2040114,-2040108,-2040102,-2040096,-2040091,-2040085,-2040079,-2040073,-2040067,-2040062,-2040056,-2040050,-2040044,-2040039,-2040033,-2040027,-2040021,-2040015,-2040010,-2040004,-2039998,-2039992,-2039987,-2039981,-2039975,-2039969,-2039963,-2039958,-2039952,-2039946,-2039940,-2039935,-2039929,-2039923,-2039917,-2039911,-2039906,-2039900,-2039894,-2039888,-2039882,-2039877,-2039871,-2039865,-2039859,-2039854,-2039848,-2039842,-2039836,-2039830,-2039825,-2039819,-2039813,-2039807,-2039801,-2039796,-2039790,-2039784,-2039778,-2039772,-2039767,-2039761,-2039755,-2039749,-2039743,-2039738,-2039732,-2039726,-2039720,-2039715,-2039709,-2039703,-2039697,-2039691,-2039686,-2039680,-2039674,-2039668,-2039662,-2039657,-2039651,-2039645,-2039639,-2039633,-2039628,-2039622,-2039616,-2039610,-2039604,-2039598,-2039593,-2039587,-2039581,-2039575,-2039569,-2039564,-2039558,-2039552,-2039546,-2039540,-2039535,-2039529,-2039523,-2039517,-2039511,-2039506,-2039500,-2039494,-2039488,-2039482,-2039476,-2039471,-2039465,-2039459,-2039453,-2039447,-2039442,-2039436,-2039430,-2039424,-2039418,-2039413,-2039407,-2039401,-2039395,-2039389,-2039383,-2039378,-2039372,-2039366,-2039360,-2039354,-2039349,-2039343,-2039337,-2039331,-2039325,-2039319,-2039314,-2039308,-2039302,-2039296,-2039290,-2039284,-2039279,-2039273,-2039267,-2039261,-2039255,-2039249,-2039244,-2039238,-2039232,-2039226,-2039220,-2039215,-2039209,-2039203,-2039197,-2039191,-2039185,-2039180,-2039174,-2039168,-2039162,-2039156,-2039150,-2039145,-2039139,-2039133,-2039127,-2039121,-2039115,-2039110,-2039104,-2039098,-2039092,-2039086,-2039080,-2039074,-2039069,-2039063,-2039057,-2039051,-2039045,-2039039,-2039034,-2039028,-2039022,-2039016,-2039010,-2039004,-2038999,-2038993,-2038987,-2038981,-2038975,-2038969,-2038963,-2038958,-2038952,-2038946,-2038940,-2038934,-2038928,-2038923,-2038917,-2038911,-2038905,-2038899,-2038893,-2038887,-2038882,-2038876,-2038870,-2038864,-2038858,-2038852,-2038846,-2038841,-2038835,-2038829,-2038823,-2038817,-2038811,-2038805,-2038800,-2038794,-2038788,-2038782,-2038776,-2038770,-2038764,-2038759,-2038753,-2038747,-2038741,-2038735,-2038729,-2038723,-2038718,-2038712,-2038706,-2038700,-2038694,-2038688,-2038682,-2038677,-2038671,-2038665,-2038659,-2038653,-2038647,-2038641,-2038635,-2038630,-2038624,-2038618,-2038612,-2038606,-2038600,-2038594,-2038589,-2038583,-2038577,-2038571,-2038565,-2038559,-2038553,-2038547,-2038542,-2038536,-2038530,-2038524,-2038518,-2038512,-2038506,-2038500,-2038495,-2038489,-2038483,-2038477,-2038471,-2038465,-2038459,-2038453,-2038448,-2038442,-2038436,-2038430,-2038424,-2038418,-2038412,-2038406,-2038400,-2038395,-2038389,-2038383,-2038377,-2038371,-2038365,-2038359,-2038353,-2038347,-2038342,-2038336,-2038330,-2038324,-2038318,-2038312,-2038306,-2038300,-2038294,-2038289,-2038283,-2038277,-2038271,-2038265,-2038259,-2038253,-2038247,-2038241,-2038236,-2038230,-2038224,-2038218,-2038212,-2038206,-2038200,-2038194,-2038188,-2038183,-2038177,-2038171,-2038165,-2038159,-2038153,-2038147,-2038141,-2038135,-2038129,-2038124,-2038118,-2038112,-2038106,-2038100,-2038094,-2038088,-2038082,-2038076,-2038070,-2038065,-2038059,-2038053,-2038047,-2038041,-2038035,-2038029,-2038023,-2038017,-2038011,-2038005,-2038000,-2037994,-2037988,-2037982,-2037976,-2037970,-2037964,-2037958,-2037952,-2037946,-2037940,-2037935,-2037929,-2037923,-2037917,-2037911,-2037905,-2037899,-2037893,-2037887,-2037881,-2037875,-2037869,-2037864,-2037858,-2037852,-2037846,-2037840,-2037834,-2037828,-2037822,-2037816,-2037810,-2037804,-2037798,-2037792,-2037787,-2037781,-2037775,-2037769,-2037763,-2037757,-2037751,-2037745,-2037739,-2037733,-2037727,-2037721,-2037715,-2037710,-2037704,-2037698,-2037692,-2037686,-2037680,-2037674,-2037668,-2037662,-2037656,-2037650,-2037644,-2037638,-2037632,-2037627,-2037621,-2037615,-2037609,-2037603,-2037597,-2037591,-2037585,-2037579,-2037573,-2037567,-2037561,-2037555,-2037549,-2037543,-2037538,-2037532,-2037526,-2037520,-2037514,-2037508,-2037502,-2037496,-2037490,-2037484,-2037478,-2037472,-2037466,-2037460,-2037454,-2037448,-2037442,-2037437,-2037431,-2037425,-2037419,-2037413,-2037407,-2037401,-2037395,-2037389,-2037383,-2037377,-2037371,-2037365,-2037359,-2037353,-2037347,-2037341,-2037335,-2037329,-2037323,-2037318,-2037312,-2037306,-2037300,-2037294,-2037288,-2037282,-2037276,-2037270,-2037264,-2037258,-2037252,-2037246,-2037240,-2037234,-2037228,-2037222,-2037216,-2037210,-2037204,-2037198,-2037192,-2037186,-2037181,-2037175,-2037169,-2037163,-2037157,-2037151,-2037145,-2037139,-2037133,-2037127,-2037121,-2037115,-2037109,-2037103,-2037097,-2037091,-2037085,-2037079,-2037073,-2037067,-2037061,-2037055,-2037049,-2037043,-2037037,-2037031,-2037025,-2037019,-2037013,-2037008,-2037002,-2036996,-2036990,-2036984,-2036978,-2036972,-2036966,-2036960,-2036954,-2036948,-2036942,-2036936,-2036930,-2036924,-2036918,-2036912,-2036906,-2036900,-2036894,-2036888,-2036882,-2036876,-2036870,-2036864,-2036858,-2036852,-2036846,-2036840,-2036834,-2036828,-2036822,-2036816,-2036810,-2036804,-2036798,-2036792,-2036786,-2036780,-2036774,-2036768,-2036762,-2036756,-2036750,-2036744,-2036738,-2036732,-2036726,-2036720,-2036714,-2036708,-2036702,-2036696,-2036690,-2036684,-2036678,-2036672,-2036666,-2036660,-2036654,-2036649,-2036643,-2036637,-2036631,-2036625,-2036619,-2036613,-2036607,-2036601,-2036595,-2036589,-2036583,-2036577,-2036571,-2036565,-2036559,-2036553,-2036547,-2036541,-2036535,-2036529,-2036523,-2036517,-2036511,-2036505,-2036499,-2036493,-2036487,-2036481,-2036474,-2036468,-2036462,-2036456,-2036450,-2036444,-2036438,-2036432,-2036426,-2036420,-2036414,-2036408,-2036402,-2036396,-2036390,-2036384,-2036378,-2036372,-2036366,-2036360,-2036354,-2036348,-2036342,-2036336,-2036330,-2036324,-2036318,-2036312,-2036306,-2036300,-2036294,-2036288,-2036282,-2036276,-2036270,-2036264,-2036258,-2036252,-2036246,-2036240,-2036234,-2036228,-2036222,-2036216,-2036210,-2036204,-2036198,-2036192,-2036186,-2036180,-2036174,-2036168,-2036162,-2036156,-2036150,-2036144,-2036138,-2036132,-2036126,-2036120,-2036113,-2036107,-2036101,-2036095,-2036089,-2036083,-2036077,-2036071,-2036065,-2036059,-2036053,-2036047,-2036041,-2036035,-2036029,-2036023,-2036017,-2036011,-2036005,-2035999,-2035993,-2035987,-2035981,-2035975,-2035969,-2035963,-2035957,-2035951,-2035945,-2035938,-2035932,-2035926,-2035920,-2035914,-2035908,-2035902,-2035896,-2035890,-2035884,-2035878,-2035872,-2035866,-2035860,-2035854,-2035848,-2035842,-2035836,-2035830,-2035824,-2035818,-2035812,-2035806,-2035799,-2035793,-2035787,-2035781,-2035775,-2035769,-2035763,-2035757,-2035751,-2035745,-2035739,-2035733,-2035727,-2035721,-2035715,-2035709,-2035703,-2035697,-2035691,-2035685,-2035678,-2035672,-2035666,-2035660,-2035654,-2035648,-2035642,-2035636,-2035630,-2035624,-2035618,-2035612,-2035606,-2035600,-2035594,-2035588,-2035582,-2035575,-2035569,-2035563,-2035557,-2035551,-2035545,-2035539,-2035533,-2035527,-2035521,-2035515,-2035509,-2035503,-2035497,-2035491,-2035484,-2035478,-2035472,-2035466,-2035460,-2035454,-2035448,-2035442,-2035436,-2035430,-2035424,-2035418,-2035412,-2035406,-2035399,-2035393,-2035387,-2035381,-2035375,-2035369,-2035363,-2035357,-2035351,-2035345,-2035339,-2035333,-2035327,-2035321,-2035314,-2035308,-2035302,-2035296,-2035290,-2035284,-2035278,-2035272,-2035266,-2035260,-2035254,-2035248,-2035241,-2035235,-2035229,-2035223,-2035217,-2035211,-2035205,-2035199,-2035193,-2035187,-2035181,-2035175,-2035168,-2035162,-2035156,-2035150,-2035144,-2035138,-2035132,-2035126,-2035120,-2035114,-2035108,-2035101,-2035095,-2035089,-2035083,-2035077,-2035071,-2035065,-2035059,-2035053,-2035047,-2035041,-2035034,-2035028,-2035022,-2035016,-2035010,-2035004,-2034998,-2034992,-2034986,-2034980,-2034973,-2034967,-2034961,-2034955,-2034949,-2034943,-2034937,-2034931,-2034925,-2034919,-2034912,-2034906,-2034900,-2034894,-2034888,-2034882,-2034876,-2034870,-2034864,-2034857,-2034851,-2034845,-2034839,-2034833,-2034827,-2034821,-2034815,-2034809,-2034803,-2034796,-2034790,-2034784,-2034778,-2034772,-2034766,-2034760,-2034754,-2034748,-2034741,-2034735,-2034729,-2034723,-2034717,-2034711,-2034705,-2034699,-2034692,-2034686,-2034680,-2034674,-2034668,-2034662,-2034656,-2034650,-2034644,-2034637,-2034631,-2034625,-2034619,-2034613,-2034607,-2034601,-2034595,-2034588,-2034582,-2034576,-2034570,-2034564,-2034558,-2034552,-2034546,-2034539,-2034533,-2034527,-2034521,-2034515,-2034509,-2034503,-2034497,-2034490,-2034484,-2034478,-2034472,-2034466,-2034460,-2034454,-2034447,-2034441,-2034435,-2034429,-2034423,-2034417,-2034411,-2034405,-2034398,-2034392,-2034386,-2034380,-2034374,-2034368,-2034362,-2034355,-2034349,-2034343,-2034337,-2034331,-2034325,-2034319,-2034312,-2034306,-2034300,-2034294,-2034288,-2034282,-2034276,-2034270,-2034263,-2034257,-2034251,-2034245,-2034239,-2034233,-2034226,-2034220,-2034214,-2034208,-2034202,-2034196,-2034190,-2034183,-2034177,-2034171,-2034165,-2034159,-2034153,-2034147,-2034140,-2034134,-2034128,-2034122,-2034116,-2034110,-2034104,-2034097,-2034091,-2034085,-2034079,-2034073,-2034067,-2034060,-2034054,-2034048,-2034042,-2034036,-2034030,-2034023,-2034017,-2034011,-2034005,-2033999,-2033993,-2033987,-2033980,-2033974,-2033968,-2033962,-2033956,-2033950,-2033943,-2033937,-2033931,-2033925,-2033919,-2033913,-2033906,-2033900,-2033894,-2033888,-2033882,-2033876,-2033869,-2033863,-2033857,-2033851,-2033845,-2033839,-2033832,-2033826,-2033820,-2033814,-2033808,-2033802,-2033795,-2033789,-2033783,-2033777,-2033771,-2033765,-2033758,-2033752,-2033746,-2033740,-2033734,-2033727,-2033721,-2033715,-2033709,-2033703,-2033697,-2033690,-2033684,-2033678,-2033672,-2033666,-2033659,-2033653,-2033647,-2033641,-2033635,-2033629,-2033622,-2033616,-2033610,-2033604,-2033598,-2033591,-2033585,-2033579,-2033573,-2033567,-2033561,-2033554,-2033548,-2033542,-2033536,-2033530,-2033523,-2033517,-2033511,-2033505,-2033499,-2033492,-2033486,-2033480,-2033474,-2033468,-2033462,-2033455,-2033449,-2033443,-2033437,-2033431,-2033424,-2033418,-2033412,-2033406,-2033400,-2033393,-2033387,-2033381,-2033375,-2033369,-2033362,-2033356,-2033350,-2033344,-2033338,-2033331,-2033325,-2033319,-2033313,-2033307,-2033300,-2033294,-2033288,-2033282,-2033276,-2033269,-2033263,-2033257,-2033251,-2033245,-2033238,-2033232,-2033226,-2033220,-2033214,-2033207,-2033201,-2033195,-2033189,-2033182,-2033176,-2033170,-2033164,-2033158,-2033151,-2033145,-2033139,-2033133,-2033127,-2033120,-2033114,-2033108,-2033102,-2033096,-2033089,-2033083,-2033077,-2033071,-2033064,-2033058,-2033052,-2033046,-2033040,-2033033,-2033027,-2033021,-2033015,-2033008,-2033002,-2032996,-2032990,-2032984,-2032977,-2032971,-2032965,-2032959,-2032952,-2032946,-2032940,-2032934,-2032928,-2032921,-2032915,-2032909,-2032903,-2032896,-2032890,-2032884,-2032878,-2032872,-2032865,-2032859,-2032853,-2032847,-2032840,-2032834,-2032828,-2032822,-2032815,-2032809,-2032803,-2032797,-2032791,-2032784,-2032778,-2032772,-2032766,-2032759,-2032753,-2032747,-2032741,-2032734,-2032728,-2032722,-2032716,-2032709,-2032703,-2032697,-2032691,-2032684,-2032678,-2032672,-2032666,-2032660,-2032653,-2032647,-2032641,-2032635,-2032628,-2032622,-2032616,-2032610,-2032603,-2032597,-2032591,-2032585,-2032578,-2032572,-2032566,-2032560,-2032553,-2032547,-2032541,-2032535,-2032528,-2032522,-2032516,-2032510,-2032503,-2032497,-2032491,-2032485,-2032478,-2032472,-2032466,-2032460,-2032453,-2032447,-2032441,-2032435,-2032428,-2032422,-2032416,-2032410,-2032403,-2032397,-2032391,-2032385,-2032378,-2032372,-2032366,-2032360,-2032353,-2032347,-2032341,-2032334,-2032328,-2032322,-2032316,-2032309,-2032303,-2032297,-2032291,-2032284,-2032278,-2032272,-2032266,-2032259,-2032253,-2032247,-2032241,-2032234,-2032228,-2032222,-2032215,-2032209,-2032203,-2032197,-2032190,-2032184,-2032178,-2032172,-2032165,-2032159,-2032153,-2032146,-2032140,-2032134,-2032128,-2032121,-2032115,-2032109,-2032103,-2032096,-2032090,-2032084,-2032077,-2032071,-2032065,-2032059,-2032052,-2032046,-2032040,-2032034,-2032027,-2032021,-2032015,-2032008,-2032002,-2031996,-2031990,-2031983,-2031977,-2031971,-2031964,-2031958,-2031952,-2031946,-2031939,-2031933,-2031927,-2031920,-2031914,-2031908,-2031902,-2031895,-2031889,-2031883,-2031876,-2031870,-2031864,-2031858,-2031851,-2031845,-2031839,-2031832,-2031826,-2031820,-2031814,-2031807,-2031801,-2031795,-2031788,-2031782,-2031776,-2031769,-2031763,-2031757,-2031751,-2031744,-2031738,-2031732,-2031725,-2031719,-2031713,-2031706,-2031700,-2031694,-2031688,-2031681,-2031675,-2031669,-2031662,-2031656,-2031650,-2031643,-2031637,-2031631,-2031625,-2031618,-2031612,-2031606,-2031599,-2031593,-2031587,-2031580,-2031574,-2031568,-2031562,-2031555,-2031549,-2031543,-2031536,-2031530,-2031524,-2031517,-2031511,-2031505,-2031498,-2031492,-2031486,-2031479,-2031473,-2031467,-2031461,-2031454,-2031448,-2031442,-2031435,-2031429,-2031423,-2031416,-2031410,-2031404,-2031397,-2031391,-2031385,-2031378,-2031372,-2031366,-2031359,-2031353,-2031347,-2031341,-2031334,-2031328,-2031322,-2031315,-2031309,-2031303,-2031296,-2031290,-2031284,-2031277,-2031271,-2031265,-2031258,-2031252,-2031246,-2031239,-2031233,-2031227,-2031220,-2031214,-2031208,-2031201,-2031195,-2031189,-2031182,-2031176,-2031170,-2031163,-2031157,-2031151,-2031144,-2031138,-2031132,-2031125,-2031119,-2031113,-2031106,-2031100,-2031094,-2031087,-2031081,-2031075,-2031068,-2031062,-2031056,-2031049,-2031043,-2031037,-2031030,-2031024,-2031018,-2031011,-2031005,-2030999,-2030992,-2030986,-2030980,-2030973,-2030967,-2030961,-2030954,-2030948,-2030942,-2030935,-2030929,-2030923,-2030916,-2030910,-2030904,-2030897,-2030891,-2030884,-2030878,-2030872,-2030865,-2030859,-2030853,-2030846,-2030840,-2030834,-2030827,-2030821,-2030815,-2030808,-2030802,-2030796,-2030789,-2030783,-2030776,-2030770,-2030764,-2030757,-2030751,-2030745,-2030738,-2030732,-2030726,-2030719,-2030713,-2030707,-2030700,-2030694,-2030687,-2030681,-2030675,-2030668,-2030662,-2030656,-2030649,-2030643,-2030637,-2030630,-2030624,-2030618,-2030611,-2030605,-2030598,-2030592,-2030586,-2030579,-2030573,-2030567,-2030560,-2030554,-2030547,-2030541,-2030535,-2030528,-2030522,-2030516,-2030509,-2030503,-2030497,-2030490,-2030484,-2030477,-2030471,-2030465,-2030458,-2030452,-2030446,-2030439,-2030433,-2030426,-2030420,-2030414,-2030407,-2030401,-2030395,-2030388,-2030382,-2030375,-2030369,-2030363,-2030356,-2030350,-2030344,-2030337,-2030331,-2030324,-2030318,-2030312,-2030305,-2030299,-2030292,-2030286,-2030280,-2030273,-2030267,-2030261,-2030254,-2030248,-2030241,-2030235,-2030229,-2030222,-2030216,-2030209,-2030203,-2030197,-2030190,-2030184,-2030178,-2030171,-2030165,-2030158,-2030152,-2030146,-2030139,-2030133,-2030126,-2030120,-2030114,-2030107,-2030101,-2030094,-2030088,-2030082,-2030075,-2030069,-2030062,-2030056,-2030050,-2030043,-2030037,-2030030,-2030024,-2030018,-2030011,-2030005,-2029998,-2029992,-2029986,-2029979,-2029973,-2029966,-2029960,-2029954,-2029947,-2029941,-2029934,-2029928,-2029922,-2029915,-2029909,-2029902,-2029896,-2029890,-2029883,-2029877,-2029870,-2029864,-2029858,-2029851,-2029845,-2029838,-2029832,-2029826,-2029819,-2029813,-2029806,-2029800,-2029793,-2029787,-2029781,-2029774,-2029768,-2029761,-2029755,-2029749,-2029742,-2029736,-2029729,-2029723,-2029716,-2029710,-2029704,-2029697,-2029691,-2029684,-2029678,-2029672,-2029665,-2029659,-2029652,-2029646,-2029639,-2029633,-2029627,-2029620,-2029614,-2029607,-2029601,-2029594,-2029588,-2029582,-2029575,-2029569,-2029562,-2029556,-2029550,-2029543,-2029537,-2029530,-2029524,-2029517,-2029511,-2029505,-2029498,-2029492,-2029485,-2029479,-2029472,-2029466,-2029460,-2029453,-2029447,-2029440,-2029434,-2029427,-2029421,-2029414,-2029408,-2029402,-2029395,-2029389,-2029382,-2029376,-2029369,-2029363,-2029357,-2029350,-2029344,-2029337,-2029331,-2029324,-2029318,-2029311,-2029305,-2029299,-2029292,-2029286,-2029279,-2029273,-2029266,-2029260,-2029253,-2029247,-2029241,-2029234,-2029228,-2029221,-2029215,-2029208,-2029202,-2029195,-2029189,-2029183,-2029176,-2029170,-2029163,-2029157,-2029150,-2029144,-2029137,-2029131,-2029125,-2029118,-2029112,-2029105,-2029099,-2029092,-2029086,-2029079,-2029073,-2029066,-2029060,-2029054,-2029047,-2029041,-2029034,-2029028,-2029021,-2029015,-2029008,-2029002,-2028995,-2028989,-2028983,-2028976,-2028970,-2028963,-2028957,-2028950,-2028944,-2028937,-2028931,-2028924,-2028918,-2028911,-2028905,-2028898,-2028892,-2028886,-2028879,-2028873,-2028866,-2028860,-2028853,-2028847,-2028840,-2028834,-2028827,-2028821,-2028814,-2028808,-2028801,-2028795,-2028789,-2028782,-2028776,-2028769,-2028763,-2028756,-2028750,-2028743,-2028737,-2028730,-2028724,-2028717,-2028711,-2028704,-2028698,-2028691,-2028685,-2028678,-2028672,-2028666,-2028659,-2028653,-2028646,-2028640,-2028633,-2028627,-2028620,-2028614,-2028607,-2028601,-2028594,-2028588,-2028581,-2028575,-2028568,-2028562,-2028555,-2028549,-2028542,-2028536,-2028529,-2028523,-2028516,-2028510,-2028503,-2028497,-2028490,-2028484,-2028477,-2028471,-2028464,-2028458,-2028452,-2028445,-2028439,-2028432,-2028426,-2028419,-2028413,-2028406,-2028400,-2028393,-2028387,-2028380,-2028374,-2028367,-2028361,-2028354,-2028348,-2028341,-2028335,-2028328,-2028322,-2028315,-2028309,-2028302,-2028296,-2028289,-2028283,-2028276,-2028270,-2028263,-2028257,-2028250,-2028244,-2028237,-2028231,-2028224,-2028218,-2028211,-2028205,-2028198,-2028192,-2028185,-2028179,-2028172,-2028166,-2028159,-2028153,-2028146,-2028140,-2028133,-2028127,-2028120,-2028113,-2028107,-2028100,-2028094,-2028087,-2028081,-2028074,-2028068,-2028061,-2028055,-2028048,-2028042,-2028035,-2028029,-2028022,-2028016,-2028009,-2028003,-2027996,-2027990,-2027983,-2027977,-2027970,-2027964,-2027957,-2027951,-2027944,-2027938,-2027931,-2027925,-2027918,-2027911,-2027905,-2027898,-2027892,-2027885,-2027879,-2027872,-2027866,-2027859,-2027853,-2027846,-2027840,-2027833,-2027827,-2027820,-2027814,-2027807,-2027801,-2027794,-2027787,-2027781,-2027774,-2027768,-2027761,-2027755,-2027748,-2027742,-2027735,-2027729,-2027722,-2027716,-2027709,-2027703,-2027696,-2027690,-2027683,-2027676,-2027670,-2027663,-2027657,-2027650,-2027644,-2027637,-2027631,-2027624,-2027618,-2027611,-2027605,-2027598,-2027591,-2027585,-2027578,-2027572,-2027565,-2027559,-2027552,-2027546,-2027539,-2027533,-2027526,-2027519,-2027513,-2027506,-2027500,-2027493,-2027487,-2027480,-2027474,-2027467,-2027461,-2027454,-2027447,-2027441,-2027434,-2027428,-2027421,-2027415,-2027408,-2027402,-2027395,-2027388,-2027382,-2027375,-2027369,-2027362,-2027356,-2027349,-2027343,-2027336,-2027330,-2027323,-2027316,-2027310,-2027303,-2027297,-2027290,-2027284,-2027277,-2027270,-2027264,-2027257,-2027251,-2027244,-2027238,-2027231,-2027225,-2027218,-2027211,-2027205,-2027198,-2027192,-2027185,-2027179,-2027172,-2027165,-2027159,-2027152,-2027146,-2027139,-2027133,-2027126,-2027120,-2027113,-2027106,-2027100,-2027093,-2027087,-2027080,-2027074,-2027067,-2027060,-2027054,-2027047,-2027041,-2027034,-2027028,-2027021,-2027014,-2027008,-2027001,-2026995,-2026988,-2026982,-2026975,-2026968,-2026962,-2026955,-2026949,-2026942,-2026935,-2026929,-2026922,-2026916,-2026909,-2026903,-2026896,-2026889,-2026883,-2026876,-2026870,-2026863,-2026857,-2026850,-2026843,-2026837,-2026830,-2026824,-2026817,-2026810,-2026804,-2026797,-2026791,-2026784,-2026777,-2026771,-2026764,-2026758,-2026751,-2026745,-2026738,-2026731,-2026725,-2026718,-2026712,-2026705,-2026698,-2026692,-2026685,-2026679,-2026672,-2026665,-2026659,-2026652,-2026646,-2026639,-2026632,-2026626,-2026619,-2026613,-2026606,-2026600,-2026593,-2026586,-2026580,-2026573,-2026567,-2026560,-2026553,-2026547,-2026540,-2026534,-2026527,-2026520,-2026514,-2026507,-2026500,-2026494,-2026487,-2026481,-2026474,-2026467,-2026461,-2026454,-2026448,-2026441,-2026434,-2026428,-2026421,-2026415,-2026408,-2026401,-2026395,-2026388,-2026382,-2026375,-2026368,-2026362,-2026355,-2026349,-2026342,-2026335,-2026329,-2026322,-2026315,-2026309,-2026302,-2026296,-2026289,-2026282,-2026276,-2026269,-2026263,-2026256,-2026249,-2026243,-2026236,-2026229,-2026223,-2026216,-2026210,-2026203,-2026196,-2026190,-2026183,-2026176,-2026170,-2026163,-2026157,-2026150,-2026143,-2026137,-2026130,-2026124,-2026117,-2026110,-2026104,-2026097,-2026090,-2026084,-2026077,-2026070,-2026064,-2026057,-2026051,-2026044,-2026037,-2026031,-2026024,-2026017,-2026011,-2026004,-2025998,-2025991,-2025984,-2025978,-2025971,-2025964,-2025958,-2025951,-2025944,-2025938,-2025931,-2025925,-2025918,-2025911,-2025905,-2025898,-2025891,-2025885,-2025878,-2025871,-2025865,-2025858,-2025852,-2025845,-2025838,-2025832,-2025825,-2025818,-2025812,-2025805,-2025798,-2025792,-2025785,-2025779,-2025772,-2025765,-2025759,-2025752,-2025745,-2025739,-2025732,-2025725,-2025719,-2025712,-2025705,-2025699,-2025692,-2025685,-2025679,-2025672,-2025666,-2025659,-2025652,-2025646,-2025639,-2025632,-2025626,-2025619,-2025612,-2025606,-2025599,-2025592,-2025586,-2025579,-2025572,-2025566,-2025559,-2025552,-2025546,-2025539,-2025532,-2025526,-2025519,-2025512,-2025506,-2025499,-2025492,-2025486,-2025479,-2025472,-2025466,-2025459,-2025452,-2025446,-2025439,-2025432,-2025426,-2025419,-2025413,-2025406,-2025399,-2025393,-2025386,-2025379,-2025373,-2025366,-2025359,-2025353,-2025346,-2025339,-2025332,-2025326,-2025319,-2025312,-2025306,-2025299,-2025292,-2025286,-2025279,-2025272,-2025266,-2025259,-2025252,-2025246,-2025239,-2025232,-2025226,-2025219,-2025212,-2025206,-2025199,-2025192,-2025186,-2025179,-2025172,-2025166,-2025159,-2025152,-2025146,-2025139,-2025132,-2025126,-2025119,-2025112,-2025106,-2025099,-2025092,-2025085,-2025079,-2025072,-2025065,-2025059,-2025052,-2025045,-2025039,-2025032,-2025025,-2025019,-2025012,-2025005,-2024999,-2024992,-2024985,-2024978,-2024972,-2024965,-2024958,-2024952,-2024945,-2024938,-2024932,-2024925,-2024918,-2024912,-2024905,-2024898,-2024891,-2024885,-2024878,-2024871,-2024865,-2024858,-2024851,-2024845,-2024838,-2024831,-2024825,-2024818,-2024811,-2024804,-2024798,-2024791,-2024784,-2024778,-2024771,-2024764,-2024758,-2024751,-2024744,-2024737,-2024731,-2024724,-2024717,-2024711,-2024704,-2024697,-2024690,-2024684,-2024677,-2024670,-2024664,-2024657,-2024650,-2024644,-2024637,-2024630,-2024623,-2024617,-2024610,-2024603,-2024597,-2024590,-2024583,-2024576,-2024570,-2024563,-2024556,-2024550,-2024543,-2024536,-2024529,-2024523,-2024516,-2024509,-2024503,-2024496,-2024489,-2024482,-2024476,-2024469,-2024462,-2024456,-2024449,-2024442,-2024435,-2024429,-2024422,-2024415,-2024409,-2024402,-2024395,-2024388,-2024382,-2024375,-2024368,-2024361,-2024355,-2024348,-2024341,-2024335,-2024328,-2024321,-2024314,-2024308,-2024301,-2024294,-2024287,-2024281,-2024274,-2024267,-2024261,-2024254,-2024247,-2024240,-2024234,-2024227,-2024220,-2024213,-2024207,-2024200,-2024193,-2024187,-2024180,-2024173,-2024166,-2024160,-2024153,-2024146,-2024139,-2024133,-2024126,-2024119,-2024112,-2024106,-2024099,-2024092,-2024085,-2024079,-2024072,-2024065,-2024058,-2024052,-2024045,-2024038,-2024032,-2024025,-2024018,-2024011,-2024005,-2023998,-2023991,-2023984,-2023978,-2023971,-2023964,-2023957,-2023951,-2023944,-2023937,-2023930,-2023924,-2023917,-2023910,-2023903,-2023897,-2023890,-2023883,-2023876,-2023870,-2023863,-2023856,-2023849,-2023843,-2023836,-2023829,-2023822,-2023816,-2023809,-2023802,-2023795,-2023789,-2023782,-2023775,-2023768,-2023762,-2023755,-2023748,-2023741,-2023734,-2023728,-2023721,-2023714,-2023707,-2023701,-2023694,-2023687,-2023680,-2023674,-2023667,-2023660,-2023653,-2023647,-2023640,-2023633,-2023626,-2023620,-2023613,-2023606,-2023599,-2023592,-2023586,-2023579,-2023572,-2023565,-2023559,-2023552,-2023545,-2023538,-2023532,-2023525,-2023518,-2023511,-2023504,-2023498,-2023491,-2023484,-2023477,-2023471,-2023464,-2023457,-2023450,-2023444,-2023437,-2023430,-2023423,-2023416,-2023410,-2023403,-2023396,-2023389,-2023383,-2023376,-2023369,-2023362,-2023355,-2023349,-2023342,-2023335,-2023328,-2023321,-2023315,-2023308,-2023301,-2023294,-2023288,-2023281,-2023274,-2023267,-2023260,-2023254,-2023247,-2023240,-2023233,-2023227,-2023220,-2023213,-2023206,-2023199,-2023193,-2023186,-2023179,-2023172,-2023165,-2023159,-2023152,-2023145,-2023138,-2023131,-2023125,-2023118,-2023111,-2023104,-2023097,-2023091,-2023084,-2023077,-2023070,-2023064,-2023057,-2023050,-2023043,-2023036,-2023030,-2023023,-2023016,-2023009,-2023002,-2022996,-2022989,-2022982,-2022975,-2022968,-2022962,-2022955,-2022948,-2022941,-2022934,-2022927,-2022921,-2022914,-2022907,-2022900,-2022893,-2022887,-2022880,-2022873,-2022866,-2022859,-2022853,-2022846,-2022839,-2022832,-2022825,-2022819,-2022812,-2022805,-2022798,-2022791,-2022785,-2022778,-2022771,-2022764,-2022757,-2022750,-2022744,-2022737,-2022730,-2022723,-2022716,-2022710,-2022703,-2022696,-2022689,-2022682,-2022675,-2022669,-2022662,-2022655,-2022648,-2022641,-2022635,-2022628,-2022621,-2022614,-2022607,-2022600,-2022594,-2022587,-2022580,-2022573,-2022566,-2022560,-2022553,-2022546,-2022539,-2022532,-2022525,-2022519,-2022512,-2022505,-2022498,-2022491,-2022484,-2022478,-2022471,-2022464,-2022457,-2022450,-2022443,-2022437,-2022430,-2022423,-2022416,-2022409,-2022402,-2022396,-2022389,-2022382,-2022375,-2022368,-2022361,-2022355,-2022348,-2022341,-2022334,-2022327,-2022320,-2022314,-2022307,-2022300,-2022293,-2022286,-2022279,-2022273,-2022266,-2022259,-2022252,-2022245,-2022238,-2022232,-2022225,-2022218,-2022211,-2022204,-2022197,-2022190,-2022184,-2022177,-2022170,-2022163,-2022156,-2022149,-2022143,-2022136,-2022129,-2022122,-2022115,-2022108,-2022101,-2022095,-2022088,-2022081,-2022074,-2022067,-2022060,-2022054,-2022047,-2022040,-2022033,-2022026,-2022019,-2022012,-2022006,-2021999,-2021992,-2021985,-2021978,-2021971,-2021964,-2021958,-2021951,-2021944,-2021937,-2021930,-2021923,-2021916,-2021910,-2021903,-2021896,-2021889,-2021882,-2021875,-2021868,-2021862,-2021855,-2021848,-2021841,-2021834,-2021827,-2021820,-2021813,-2021807,-2021800,-2021793,-2021786,-2021779,-2021772,-2021765,-2021759,-2021752,-2021745,-2021738,-2021731,-2021724,-2021717,-2021710,-2021704,-2021697,-2021690,-2021683,-2021676,-2021669,-2021662,-2021655,-2021649,-2021642,-2021635,-2021628,-2021621,-2021614,-2021607,-2021600,-2021594,-2021587,-2021580,-2021573,-2021566,-2021559,-2021552,-2021545,-2021539,-2021532,-2021525,-2021518,-2021511,-2021504,-2021497,-2021490,-2021484,-2021477,-2021470,-2021463,-2021456,-2021449,-2021442,-2021435,-2021428,-2021422,-2021415,-2021408,-2021401,-2021394,-2021387,-2021380,-2021373,-2021366,-2021360,-2021353,-2021346,-2021339,-2021332,-2021325,-2021318,-2021311,-2021304,-2021298,-2021291,-2021284,-2021277,-2021270,-2021263,-2021256,-2021249,-2021242,-2021235,-2021229,-2021222,-2021215,-2021208,-2021201,-2021194,-2021187,-2021180,-2021173,-2021166,-2021160,-2021153,-2021146,-2021139,-2021132,-2021125,-2021118,-2021111,-2021104,-2021097,-2021091,-2021084,-2021077,-2021070,-2021063,-2021056,-2021049,-2021042,-2021035,-2021028,-2021021,-2021015,-2021008,-2021001,-2020994,-2020987,-2020980,-2020973,-2020966,-2020959,-2020952,-2020945,-2020939,-2020932,-2020925,-2020918,-2020911,-2020904,-2020897,-2020890,-2020883,-2020876,-2020869,-2020863,-2020856,-2020849,-2020842,-2020835,-2020828,-2020821,-2020814,-2020807,-2020800,-2020793,-2020786,-2020779,-2020773,-2020766,-2020759,-2020752,-2020745,-2020738,-2020731,-2020724,-2020717,-2020710,-2020703,-2020696,-2020689,-2020683,-2020676,-2020669,-2020662,-2020655,-2020648,-2020641,-2020634,-2020627,-2020620,-2020613,-2020606,-2020599,-2020592,-2020586,-2020579,-2020572,-2020565,-2020558,-2020551,-2020544,-2020537,-2020530,-2020523,-2020516,-2020509,-2020502,-2020495,-2020488,-2020482,-2020475,-2020468,-2020461,-2020454,-2020447,-2020440,-2020433,-2020426,-2020419,-2020412,-2020405,-2020398,-2020391,-2020384,-2020377,-2020370,-2020364,-2020357,-2020350,-2020343,-2020336,-2020329,-2020322,-2020315,-2020308,-2020301,-2020294,-2020287,-2020280,-2020273,-2020266,-2020259,-2020252,-2020245,-2020238,-2020232,-2020225,-2020218,-2020211,-2020204,-2020197,-2020190,-2020183,-2020176,-2020169,-2020162,-2020155,-2020148,-2020141,-2020134,-2020127,-2020120,-2020113,-2020106,-2020099,-2020092,-2020085,-2020078,-2020072,-2020065,-2020058,-2020051,-2020044,-2020037,-2020030,-2020023,-2020016,-2020009,-2020002,-2019995,-2019988,-2019981,-2019974,-2019967,-2019960,-2019953,-2019946,-2019939,-2019932,-2019925,-2019918,-2019911,-2019904,-2019897,-2019890,-2019883,-2019877,-2019870,-2019863,-2019856,-2019849,-2019842,-2019835,-2019828,-2019821,-2019814,-2019807,-2019800,-2019793,-2019786,-2019779,-2019772,-2019765,-2019758,-2019751,-2019744,-2019737,-2019730,-2019723,-2019716,-2019709,-2019702,-2019695,-2019688,-2019681,-2019674,-2019667,-2019660,-2019653,-2019646,-2019639,-2019632,-2019625,-2019618,-2019611,-2019604,-2019597,-2019590,-2019583,-2019576,-2019569,-2019562,-2019555,-2019548,-2019541,-2019535,-2019528,-2019521,-2019514,-2019507,-2019500,-2019493,-2019486,-2019479,-2019472,-2019465,-2019458,-2019451,-2019444,-2019437,-2019430,-2019423,-2019416,-2019409,-2019402,-2019395,-2019388,-2019381,-2019374,-2019367,-2019360,-2019353,-2019346,-2019339,-2019332,-2019325,-2019318,-2019311,-2019304,-2019297,-2019290,-2019283,-2019276,-2019269,-2019262,-2019255,-2019248,-2019241,-2019234,-2019227,-2019220,-2019213,-2019206,-2019199,-2019192,-2019185,-2019178,-2019171,-2019164,-2019157,-2019150,-2019143,-2019136,-2019129,-2019122,-2019115,-2019107,-2019100,-2019093,-2019086,-2019079,-2019072,-2019065,-2019058,-2019051,-2019044,-2019037,-2019030,-2019023,-2019016,-2019009,-2019002,-2018995,-2018988,-2018981,-2018974,-2018967,-2018960,-2018953,-2018946,-2018939,-2018932,-2018925,-2018918,-2018911,-2018904,-2018897,-2018890,-2018883,-2018876,-2018869,-2018862,-2018855,-2018848,-2018841,-2018834,-2018827,-2018820,-2018813,-2018806,-2018799,-2018792,-2018785,-2018778,-2018771,-2018763,-2018756,-2018749,-2018742,-2018735,-2018728,-2018721,-2018714,-2018707,-2018700,-2018693,-2018686,-2018679,-2018672,-2018665,-2018658,-2018651,-2018644,-2018637,-2018630,-2018623,-2018616,-2018609,-2018602,-2018595,-2018588,-2018581,-2018574,-2018566,-2018559,-2018552,-2018545,-2018538,-2018531,-2018524,-2018517,-2018510,-2018503,-2018496,-2018489,-2018482,-2018475,-2018468,-2018461,-2018454,-2018447,-2018440,-2018433,-2018426,-2018419,-2018412,-2018404,-2018397,-2018390,-2018383,-2018376,-2018369,-2018362,-2018355,-2018348,-2018341,-2018334,-2018327,-2018320,-2018313,-2018306,-2018299,-2018292,-2018285,-2018278,-2018270,-2018263,-2018256,-2018249,-2018242,-2018235,-2018228,-2018221,-2018214,-2018207,-2018200,-2018193,-2018186,-2018179,-2018172,-2018165,-2018158,-2018150,-2018143,-2018136,-2018129,-2018122,-2018115,-2018108,-2018101,-2018094,-2018087,-2018080,-2018073,-2018066,-2018059,-2018052,-2018044,-2018037,-2018030,-2018023,-2018016,-2018009,-2018002,-2017995,-2017988,-2017981,-2017974,-2017967,-2017960,-2017953,-2017945,-2017938,-2017931,-2017924,-2017917,-2017910,-2017903,-2017896,-2017889,-2017882,-2017875,-2017868,-2017861,-2017853,-2017846,-2017839,-2017832,-2017825,-2017818,-2017811,-2017804,-2017797,-2017790,-2017783,-2017776,-2017769,-2017761,-2017754,-2017747,-2017740,-2017733,-2017726,-2017719,-2017712,-2017705,-2017698,-2017691,-2017683,-2017676,-2017669,-2017662,-2017655,-2017648,-2017641,-2017634,-2017627,-2017620,-2017613,-2017606,-2017598,-2017591,-2017584,-2017577,-2017570,-2017563,-2017556,-2017549,-2017542,-2017535,-2017527,-2017520,-2017513,-2017506,-2017499,-2017492,-2017485,-2017478,-2017471,-2017464,-2017456,-2017449,-2017442,-2017435,-2017428,-2017421,-2017414,-2017407,-2017400,-2017393,-2017385,-2017378,-2017371,-2017364,-2017357,-2017350,-2017343,-2017336,-2017329,-2017322,-2017314,-2017307,-2017300,-2017293,-2017286,-2017279,-2017272,-2017265,-2017258,-2017250,-2017243,-2017236,-2017229,-2017222,-2017215,-2017208,-2017201,-2017194,-2017186,-2017179,-2017172,-2017165,-2017158,-2017151,-2017144,-2017137,-2017130,-2017122,-2017115,-2017108,-2017101,-2017094,-2017087,-2017080,-2017073,-2017065,-2017058,-2017051,-2017044,-2017037,-2017030,-2017023,-2017016,-2017008,-2017001,-2016994,-2016987,-2016980,-2016973,-2016966,-2016959,-2016951,-2016944,-2016937,-2016930,-2016923,-2016916,-2016909,-2016902,-2016894,-2016887,-2016880,-2016873,-2016866,-2016859,-2016852,-2016845,-2016837,-2016830,-2016823,-2016816,-2016809,-2016802,-2016795,-2016787,-2016780,-2016773,-2016766,-2016759,-2016752,-2016745,-2016738,-2016730,-2016723,-2016716,-2016709,-2016702,-2016695,-2016688,-2016680,-2016673,-2016666,-2016659,-2016652,-2016645,-2016638,-2016630,-2016623,-2016616,-2016609,-2016602,-2016595,-2016588,-2016580,-2016573,-2016566,-2016559,-2016552,-2016545,-2016538,-2016530,-2016523,-2016516,-2016509,-2016502,-2016495,-2016488,-2016480,-2016473,-2016466,-2016459,-2016452,-2016445,-2016437,-2016430,-2016423,-2016416,-2016409,-2016402,-2016395,-2016387,-2016380,-2016373,-2016366,-2016359,-2016352,-2016344,-2016337,-2016330,-2016323,-2016316,-2016309,-2016301,-2016294,-2016287,-2016280,-2016273,-2016266,-2016258,-2016251,-2016244,-2016237,-2016230,-2016223,-2016216,-2016208,-2016201,-2016194,-2016187,-2016180,-2016173,-2016165,-2016158,-2016151,-2016144,-2016137,-2016130,-2016122,-2016115,-2016108,-2016101,-2016094,-2016086,-2016079,-2016072,-2016065,-2016058,-2016051,-2016043,-2016036,-2016029,-2016022,-2016015,-2016008,-2016000,-2015993,-2015986,-2015979,-2015972,-2015965,-2015957,-2015950,-2015943,-2015936,-2015929,-2015921,-2015914,-2015907,-2015900,-2015893,-2015886,-2015878,-2015871,-2015864,-2015857,-2015850,-2015842,-2015835,-2015828,-2015821,-2015814,-2015807,-2015799,-2015792,-2015785,-2015778,-2015771,-2015763,-2015756,-2015749,-2015742,-2015735,-2015727,-2015720,-2015713,-2015706,-2015699,-2015691,-2015684,-2015677,-2015670,-2015663,-2015656,-2015648,-2015641,-2015634,-2015627,-2015620,-2015612,-2015605,-2015598,-2015591,-2015584,-2015576,-2015569,-2015562,-2015555,-2015548,-2015540,-2015533,-2015526,-2015519,-2015512,-2015504,-2015497,-2015490,-2015483,-2015476,-2015468,-2015461,-2015454,-2015447,-2015440,-2015432,-2015425,-2015418,-2015411,-2015404,-2015396,-2015389,-2015382,-2015375,-2015367,-2015360,-2015353,-2015346,-2015339,-2015331,-2015324,-2015317,-2015310,-2015303,-2015295,-2015288,-2015281,-2015274,-2015267,-2015259,-2015252,-2015245,-2015238,-2015230,-2015223,-2015216,-2015209,-2015202,-2015194,-2015187,-2015180,-2015173,-2015165,-2015158,-2015151,-2015144,-2015137,-2015129,-2015122,-2015115,-2015108,-2015100,-2015093,-2015086,-2015079,-2015072,-2015064,-2015057,-2015050,-2015043,-2015035,-2015028,-2015021,-2015014,-2015007,-2014999,-2014992,-2014985,-2014978,-2014970,-2014963,-2014956,-2014949,-2014941,-2014934,-2014927,-2014920,-2014913,-2014905,-2014898,-2014891,-2014884,-2014876,-2014869,-2014862,-2014855,-2014847,-2014840,-2014833,-2014826,-2014819,-2014811,-2014804,-2014797,-2014790,-2014782,-2014775,-2014768,-2014761,-2014753,-2014746,-2014739,-2014732,-2014724,-2014717,-2014710,-2014703,-2014695,-2014688,-2014681,-2014674,-2014666,-2014659,-2014652,-2014645,-2014637,-2014630,-2014623,-2014616,-2014608,-2014601,-2014594,-2014587,-2014579,-2014572,-2014565,-2014558,-2014550,-2014543,-2014536,-2014529,-2014521,-2014514,-2014507,-2014500,-2014492,-2014485,-2014478,-2014471,-2014463,-2014456,-2014449,-2014442,-2014434,-2014427,-2014420,-2014413,-2014405,-2014398,-2014391,-2014384,-2014376,-2014369,-2014362,-2014355,-2014347,-2014340,-2014333,-2014325,-2014318,-2014311,-2014304,-2014296,-2014289,-2014282,-2014275,-2014267,-2014260,-2014253,-2014246,-2014238,-2014231,-2014224,-2014217,-2014209,-2014202,-2014195,-2014187,-2014180,-2014173,-2014166,-2014158,-2014151,-2014144,-2014137,-2014129,-2014122,-2014115,-2014107,-2014100,-2014093,-2014086,-2014078,-2014071,-2014064,-2014057,-2014049,-2014042,-2014035,-2014027,-2014020,-2014013,-2014006,-2013998,-2013991,-2013984,-2013976,-2013969,-2013962,-2013955,-2013947,-2013940,-2013933,-2013925,-2013918,-2013911,-2013904,-2013896,-2013889,-2013882,-2013874,-2013867,-2013860,-2013853,-2013845,-2013838,-2013831,-2013823,-2013816,-2013809,-2013802,-2013794,-2013787,-2013780,-2013772,-2013765,-2013758,-2013751,-2013743,-2013736,-2013729,-2013721,-2013714,-2013707,-2013700,-2013692,-2013685,-2013678,-2013670,-2013663,-2013656,-2013648,-2013641,-2013634,-2013627,-2013619,-2013612,-2013605,-2013597,-2013590,-2013583,-2013575,-2013568,-2013561,-2013554,-2013546,-2013539,-2013532,-2013524,-2013517,-2013510,-2013502,-2013495,-2013488,-2013480,-2013473,-2013466,-2013459,-2013451,-2013444,-2013437,-2013429,-2013422,-2013415,-2013407,-2013400,-2013393,-2013385,-2013378,-2013371,-2013364,-2013356,-2013349,-2013342,-2013334,-2013327,-2013320,-2013312,-2013305,-2013298,-2013290,-2013283,-2013276,-2013268,-2013261,-2013254,-2013246,-2013239,-2013232,-2013225,-2013217,-2013210,-2013203,-2013195,-2013188,-2013181,-2013173,-2013166,-2013159,-2013151,-2013144,-2013137,-2013129,-2013122,-2013115,-2013107,-2013100,-2013093,-2013085,-2013078,-2013071,-2013063,-2013056,-2013049,-2013041,-2013034,-2013027,-2013019,-2013012,-2013005,-2012997,-2012990,-2012983,-2012975,-2012968,-2012961,-2012953,-2012946,-2012939,-2012931,-2012924,-2012917,-2012909,-2012902,-2012895,-2012887,-2012880,-2012873,-2012865,-2012858,-2012851,-2012843,-2012836,-2012829,-2012821,-2012814,-2012807,-2012799,-2012792,-2012785,-2012777,-2012770,-2012763,-2012755,-2012748,-2012741,-2012733,-2012726,-2012719,-2012711,-2012704,-2012697,-2012689,-2012682,-2012675,-2012667,-2012660,-2012652,-2012645,-2012638,-2012630,-2012623,-2012616,-2012608,-2012601,-2012594,-2012586,-2012579,-2012572,-2012564,-2012557,-2012550,-2012542,-2012535,-2012528,-2012520,-2012513,-2012505,-2012498,-2012491,-2012483,-2012476,-2012469,-2012461,-2012454,-2012447,-2012439,-2012432,-2012424,-2012417,-2012410,-2012402,-2012395,-2012388,-2012380,-2012373,-2012366,-2012358,-2012351,-2012344,-2012336,-2012329,-2012321,-2012314,-2012307,-2012299,-2012292,-2012285,-2012277,-2012270,-2012262,-2012255,-2012248,-2012240,-2012233,-2012226,-2012218,-2012211,-2012204,-2012196,-2012189,-2012181,-2012174,-2012167,-2012159,-2012152,-2012145,-2012137,-2012130,-2012122,-2012115,-2012108,-2012100,-2012093,-2012086,-2012078,-2012071,-2012063,-2012056,-2012049,-2012041,-2012034,-2012027,-2012019,-2012012,-2012004,-2011997,-2011990,-2011982,-2011975,-2011967,-2011960,-2011953,-2011945,-2011938,-2011931,-2011923,-2011916,-2011908,-2011901,-2011894,-2011886,-2011879,-2011871,-2011864,-2011857,-2011849,-2011842,-2011834,-2011827,-2011820,-2011812,-2011805,-2011798,-2011790,-2011783,-2011775,-2011768,-2011761,-2011753,-2011746,-2011738,-2011731,-2011724,-2011716,-2011709,-2011701,-2011694,-2011687,-2011679,-2011672,-2011664,-2011657,-2011650,-2011642,-2011635,-2011627,-2011620,-2011613,-2011605,-2011598,-2011590,-2011583,-2011576,-2011568,-2011561,-2011553,-2011546,-2011539,-2011531,-2011524,-2011516,-2011509,-2011502,-2011494,-2011487,-2011479,-2011472,-2011465,-2011457,-2011450,-2011442,-2011435,-2011427,-2011420,-2011413,-2011405,-2011398,-2011390,-2011383,-2011376,-2011368,-2011361,-2011353,-2011346,-2011339,-2011331,-2011324,-2011316,-2011309,-2011301,-2011294,-2011287,-2011279,-2011272,-2011264,-2011257,-2011250,-2011242,-2011235,-2011227,-2011220,-2011212,-2011205,-2011198,-2011190,-2011183,-2011175,-2011168,-2011160,-2011153,-2011146,-2011138,-2011131,-2011123,-2011116,-2011108,-2011101,-2011094,-2011086,-2011079,-2011071,-2011064,-2011056,-2011049,-2011042,-2011034,-2011027,-2011019,-2011012,-2011004,-2010997,-2010990,-2010982,-2010975,-2010967,-2010960,-2010952,-2010945,-2010938,-2010930,-2010923,-2010915,-2010908,-2010900,-2010893,-2010885,-2010878,-2010871,-2010863,-2010856,-2010848,-2010841,-2010833,-2010826,-2010819,-2010811,-2010804,-2010796,-2010789,-2010781,-2010774,-2010766,-2010759,-2010752,-2010744,-2010737,-2010729,-2010722,-2010714,-2010707,-2010699,-2010692,-2010685,-2010677,-2010670,-2010662,-2010655,-2010647,-2010640,-2010632,-2010625,-2010617,-2010610,-2010603,-2010595,-2010588,-2010580,-2010573,-2010565,-2010558,-2010550,-2010543,-2010535,-2010528,-2010521,-2010513,-2010506,-2010498,-2010491,-2010483,-2010476,-2010468,-2010461,-2010453,-2010446,-2010439,-2010431,-2010424,-2010416,-2010409,-2010401,-2010394,-2010386,-2010379,-2010371,-2010364,-2010356,-2010349,-2010342,-2010334,-2010327,-2010319,-2010312,-2010304,-2010297,-2010289,-2010282,-2010274,-2010267,-2010259,-2010252,-2010244,-2010237,-2010229,-2010222,-2010215,-2010207,-2010200,-2010192,-2010185,-2010177,-2010170,-2010162,-2010155,-2010147,-2010140,-2010132,-2010125,-2010117,-2010110,-2010102,-2010095,-2010087,-2010080,-2010073,-2010065,-2010058,-2010050,-2010043,-2010035,-2010028,-2010020,-2010013,-2010005,-2009998,-2009990,-2009983,-2009975,-2009968,-2009960,-2009953,-2009945,-2009938,-2009930,-2009923,-2009915,-2009908,-2009900,-2009893,-2009885,-2009878,-2009870,-2009863,-2009855,-2009848,-2009841,-2009833,-2009826,-2009818,-2009811,-2009803,-2009796,-2009788,-2009781,-2009773,-2009766,-2009758,-2009751,-2009743,-2009736,-2009728,-2009721,-2009713,-2009706,-2009698,-2009691,-2009683,-2009676,-2009668,-2009661,-2009653,-2009646,-2009638,-2009631,-2009623,-2009616,-2009608,-2009601,-2009593,-2009586,-2009578,-2009571,-2009563,-2009556,-2009548,-2009541,-2009533,-2009526,-2009518,-2009511,-2009503,-2009496,-2009488,-2009481,-2009473,-2009466,-2009458,-2009451,-2009443,-2009435,-2009428,-2009420,-2009413,-2009405,-2009398,-2009390,-2009383,-2009375,-2009368,-2009360,-2009353,-2009345,-2009338,-2009330,-2009323,-2009315,-2009308,-2009300,-2009293,-2009285,-2009278,-2009270,-2009263,-2009255,-2009248,-2009240,-2009233,-2009225,-2009218,-2009210,-2009202,-2009195,-2009187,-2009180,-2009172,-2009165,-2009157,-2009150,-2009142,-2009135,-2009127,-2009120,-2009112,-2009105,-2009097,-2009090,-2009082,-2009075,-2009067,-2009059,-2009052,-2009044,-2009037,-2009029,-2009022,-2009014,-2009007,-2008999,-2008992,-2008984,-2008977,-2008969,-2008962,-2008954,-2008947,-2008939,-2008931,-2008924,-2008916,-2008909,-2008901,-2008894,-2008886,-2008879,-2008871,-2008864,-2008856,-2008849,-2008841,-2008833,-2008826,-2008818,-2008811,-2008803,-2008796,-2008788,-2008781,-2008773,-2008766,-2008758,-2008750,-2008743,-2008735,-2008728,-2008720,-2008713,-2008705,-2008698,-2008690,-2008683,-2008675,-2008667,-2008660,-2008652,-2008645,-2008637,-2008630,-2008622,-2008615,-2008607,-2008600,-2008592,-2008584,-2008577,-2008569,-2008562,-2008554,-2008547,-2008539,-2008532,-2008524,-2008516,-2008509,-2008501,-2008494,-2008486,-2008479,-2008471,-2008464,-2008456,-2008448,-2008441,-2008433,-2008426,-2008418,-2008411,-2008403,-2008395,-2008388,-2008380,-2008373,-2008365,-2008358,-2008350,-2008343,-2008335,-2008327,-2008320,-2008312,-2008305,-2008297,-2008290,-2008282,-2008274,-2008267,-2008259,-2008252,-2008244,-2008237,-2008229,-2008221,-2008214,-2008206,-2008199,-2008191,-2008184,-2008176,-2008168,-2008161,-2008153,-2008146,-2008138,-2008131,-2008123,-2008115,-2008108,-2008100,-2008093,-2008085,-2008078,-2008070,-2008062,-2008055,-2008047,-2008040,-2008032,-2008024,-2008017,-2008009,-2008002,-2007994,-2007987,-2007979,-2007971,-2007964,-2007956,-2007949,-2007941,-2007933,-2007926,-2007918,-2007911,-2007903,-2007896,-2007888,-2007880,-2007873,-2007865,-2007858,-2007850,-2007842,-2007835,-2007827,-2007820,-2007812,-2007805,-2007797,-2007789,-2007782,-2007774,-2007767,-2007759,-2007751,-2007744,-2007736,-2007729,-2007721,-2007713,-2007706,-2007698,-2007691,-2007683,-2007675,-2007668,-2007660,-2007653,-2007645,-2007637,-2007630,-2007622,-2007615,-2007607,-2007599,-2007592,-2007584,-2007577,-2007569,-2007561,-2007554,-2007546,-2007539,-2007531,-2007523,-2007516,-2007508,-2007501,-2007493,-2007485,-2007478,-2007470,-2007463,-2007455,-2007447,-2007440,-2007432,-2007424,-2007417,-2007409,-2007402,-2007394,-2007386,-2007379,-2007371,-2007364,-2007356,-2007348,-2007341,-2007333,-2007326,-2007318,-2007310,-2007303,-2007295,-2007287,-2007280,-2007272,-2007265,-2007257,-2007249,-2007242,-2007234,-2007226,-2007219,-2007211,-2007204,-2007196,-2007188,-2007181,-2007173,-2007166,-2007158,-2007150,-2007143,-2007135,-2007127,-2007120,-2007112,-2007105,-2007097,-2007089,-2007082,-2007074,-2007066,-2007059,-2007051,-2007044,-2007036,-2007028,-2007021,-2007013,-2007005,-2006998,-2006990,-2006982,-2006975,-2006967,-2006960,-2006952,-2006944,-2006937,-2006929,-2006921,-2006914,-2006906,-2006899,-2006891,-2006883,-2006876,-2006868,-2006860,-2006853,-2006845,-2006837,-2006830,-2006822,-2006814,-2006807,-2006799,-2006792,-2006784,-2006776,-2006769,-2006761,-2006753,-2006746,-2006738,-2006730,-2006723,-2006715,-2006708,-2006700,-2006692,-2006685,-2006677,-2006669,-2006662,-2006654,-2006646,-2006639,-2006631,-2006623,-2006616,-2006608,-2006600,-2006593,-2006585,-2006577,-2006570,-2006562,-2006555,-2006547,-2006539,-2006532,-2006524,-2006516,-2006509,-2006501,-2006493,-2006486,-2006478,-2006470,-2006463,-2006455,-2006447,-2006440,-2006432,-2006424,-2006417,-2006409,-2006401,-2006394,-2006386,-2006378,-2006371,-2006363,-2006355,-2006348,-2006340,-2006332,-2006325,-2006317,-2006309,-2006302,-2006294,-2006286,-2006279,-2006271,-2006263,-2006256,-2006248,-2006240,-2006233,-2006225,-2006217,-2006210,-2006202,-2006194,-2006187,-2006179,-2006171,-2006164,-2006156,-2006148,-2006141,-2006133,-2006125,-2006118,-2006110,-2006102,-2006095,-2006087,-2006079,-2006072,-2006064,-2006056,-2006049,-2006041,-2006033,-2006026,-2006018,-2006010,-2006003,-2005995,-2005987,-2005980,-2005972,-2005964,-2005957,-2005949,-2005941,-2005933,-2005926,-2005918,-2005910,-2005903,-2005895,-2005887,-2005880,-2005872,-2005864,-2005857,-2005849,-2005841,-2005834,-2005826,-2005818,-2005811,-2005803,-2005795,-2005787,-2005780,-2005772,-2005764,-2005757,-2005749,-2005741,-2005734,-2005726,-2005718,-2005711,-2005703,-2005695,-2005687,-2005680,-2005672,-2005664,-2005657,-2005649,-2005641,-2005634,-2005626,-2005618,-2005610,-2005603,-2005595,-2005587,-2005580,-2005572,-2005564,-2005557,-2005549,-2005541,-2005533,-2005526,-2005518,-2005510,-2005503,-2005495,-2005487,-2005480,-2005472,-2005464,-2005456,-2005449,-2005441,-2005433,-2005426,-2005418,-2005410,-2005402,-2005395,-2005387,-2005379,-2005372,-2005364,-2005356,-2005349,-2005341,-2005333,-2005325,-2005318,-2005310,-2005302,-2005295,-2005287,-2005279,-2005271,-2005264,-2005256,-2005248,-2005241,-2005233,-2005225,-2005217,-2005210,-2005202,-2005194,-2005187,-2005179,-2005171,-2005163,-2005156,-2005148,-2005140,-2005132,-2005125,-2005117,-2005109,-2005102,-2005094,-2005086,-2005078,-2005071,-2005063,-2005055,-2005048,-2005040,-2005032,-2005024,-2005017,-2005009,-2005001,-2004993,-2004986,-2004978,-2004970,-2004963,-2004955,-2004947,-2004939,-2004932,-2004924,-2004916,-2004908,-2004901,-2004893,-2004885,-2004877,-2004870,-2004862,-2004854,-2004847,-2004839,-2004831,-2004823,-2004816,-2004808,-2004800,-2004792,-2004785,-2004777,-2004769,-2004761,-2004754,-2004746,-2004738,-2004730,-2004723,-2004715,-2004707,-2004699,-2004692,-2004684,-2004676,-2004669,-2004661,-2004653,-2004645,-2004638,-2004630,-2004622,-2004614,-2004607,-2004599,-2004591,-2004583,-2004576,-2004568,-2004560,-2004552,-2004545,-2004537,-2004529,-2004521,-2004514,-2004506,-2004498,-2004490,-2004483,-2004475,-2004467,-2004459,-2004452,-2004444,-2004436,-2004428,-2004421,-2004413,-2004405,-2004397,-2004389,-2004382,-2004374,-2004366,-2004358,-2004351,-2004343,-2004335,-2004327,-2004320,-2004312,-2004304,-2004296,-2004289,-2004281,-2004273,-2004265,-2004258,-2004250,-2004242,-2004234,-2004227,-2004219,-2004211,-2004203,-2004195,-2004188,-2004180,-2004172,-2004164,-2004157,-2004149,-2004141,-2004133,-2004126,-2004118,-2004110,-2004102,-2004094,-2004087,-2004079,-2004071,-2004063,-2004056,-2004048,-2004040,-2004032,-2004025,-2004017,-2004009,-2004001,-2003993,-2003986,-2003978,-2003970,-2003962,-2003955,-2003947,-2003939,-2003931,-2003923,-2003916,-2003908,-2003900,-2003892,-2003884,-2003877,-2003869,-2003861,-2003853,-2003846,-2003838,-2003830,-2003822,-2003814,-2003807,-2003799,-2003791,-2003783,-2003776,-2003768,-2003760,-2003752,-2003744,-2003737,-2003729,-2003721,-2003713,-2003705,-2003698,-2003690,-2003682,-2003674,-2003666,-2003659,-2003651,-2003643,-2003635,-2003628,-2003620,-2003612,-2003604,-2003596,-2003589,-2003581,-2003573,-2003565,-2003557,-2003550,-2003542,-2003534,-2003526,-2003518,-2003511,-2003503,-2003495,-2003487,-2003479,-2003472,-2003464,-2003456,-2003448,-2003440,-2003433,-2003425,-2003417,-2003409,-2003401,-2003394,-2003386,-2003378,-2003370,-2003362,-2003355,-2003347,-2003339,-2003331,-2003323,-2003315,-2003308,-2003300,-2003292,-2003284,-2003276,-2003269,-2003261,-2003253,-2003245,-2003237,-2003230,-2003222,-2003214,-2003206,-2003198,-2003190,-2003183,-2003175,-2003167,-2003159,-2003151,-2003144,-2003136,-2003128,-2003120,-2003112,-2003104,-2003097,-2003089,-2003081,-2003073,-2003065,-2003058,-2003050,-2003042,-2003034,-2003026,-2003018,-2003011,-2003003,-2002995,-2002987,-2002979,-2002972,-2002964,-2002956,-2002948,-2002940,-2002932,-2002925,-2002917,-2002909,-2002901,-2002893,-2002885,-2002878,-2002870,-2002862,-2002854,-2002846,-2002838,-2002831,-2002823,-2002815,-2002807,-2002799,-2002791,-2002784,-2002776,-2002768,-2002760,-2002752,-2002744,-2002737,-2002729,-2002721,-2002713,-2002705,-2002697,-2002690,-2002682,-2002674,-2002666,-2002658,-2002650,-2002643,-2002635,-2002627,-2002619,-2002611,-2002603,-2002596,-2002588,-2002580,-2002572,-2002564,-2002556,-2002548,-2002541,-2002533,-2002525,-2002517,-2002509,-2002501,-2002494,-2002486,-2002478,-2002470,-2002462,-2002454,-2002446,-2002439,-2002431,-2002423,-2002415,-2002407,-2002399,-2002391,-2002384,-2002376,-2002368,-2002360,-2002352,-2002344,-2002336,-2002329,-2002321,-2002313,-2002305,-2002297,-2002289,-2002281,-2002274,-2002266,-2002258,-2002250,-2002242,-2002234,-2002226,-2002219,-2002211,-2002203,-2002195,-2002187,-2002179,-2002171,-2002164,-2002156,-2002148,-2002140,-2002132,-2002124,-2002116,-2002109,-2002101,-2002093,-2002085,-2002077,-2002069,-2002061,-2002053,-2002046,-2002038,-2002030,-2002022,-2002014,-2002006,-2001998,-2001991,-2001983,-2001975,-2001967,-2001959,-2001951,-2001943,-2001935,-2001928,-2001920,-2001912,-2001904,-2001896,-2001888,-2001880,-2001872,-2001865,-2001857,-2001849,-2001841,-2001833,-2001825,-2001817,-2001809,-2001801,-2001794,-2001786,-2001778,-2001770,-2001762,-2001754,-2001746,-2001738,-2001731,-2001723,-2001715,-2001707,-2001699,-2001691,-2001683,-2001675,-2001667,-2001660,-2001652,-2001644,-2001636,-2001628,-2001620,-2001612,-2001604,-2001596,-2001589,-2001581,-2001573,-2001565,-2001557,-2001549,-2001541,-2001533,-2001525,-2001518,-2001510,-2001502,-2001494,-2001486,-2001478,-2001470,-2001462,-2001454,-2001446,-2001439,-2001431,-2001423,-2001415,-2001407,-2001399,-2001391,-2001383,-2001375,-2001367,-2001360,-2001352,-2001344,-2001336,-2001328,-2001320,-2001312,-2001304,-2001296,-2001288,-2001281,-2001273,-2001265,-2001257,-2001249,-2001241,-2001233,-2001225,-2001217,-2001209,-2001201,-2001194,-2001186,-2001178,-2001170,-2001162,-2001154,-2001146,-2001138,-2001130,-2001122,-2001114,-2001107,-2001099,-2001091,-2001083,-2001075,-2001067,-2001059,-2001051,-2001043,-2001035,-2001027,-2001019,-2001012,-2001004,-2000996,-2000988,-2000980,-2000972,-2000964,-2000956,-2000948,-2000940,-2000932,-2000924,-2000917,-2000909,-2000901,-2000893,-2000885,-2000877,-2000869,-2000861,-2000853,-2000845,-2000837,-2000829,-2000821,-2000814,-2000806,-2000798,-2000790,-2000782,-2000774,-2000766,-2000758,-2000750,-2000742,-2000734,-2000726,-2000718,-2000710,-2000703,-2000695,-2000687,-2000679,-2000671,-2000663,-2000655,-2000647,-2000639,-2000631,-2000623,-2000615,-2000607,-2000599,-2000591,-2000583,-2000576,-2000568,-2000560,-2000552,-2000544,-2000536,-2000528,-2000520,-2000512,-2000504,-2000496,-2000488,-2000480,-2000472,-2000464,-2000456,-2000448,-2000441,-2000433,-2000425,-2000417,-2000409,-2000401,-2000393,-2000385,-2000377,-2000369,-2000361,-2000353,-2000345,-2000337,-2000329,-2000321,-2000313,-2000305,-2000297,-2000290,-2000282,-2000274,-2000266,-2000258,-2000250,-2000242,-2000234,-2000226,-2000218,-2000210,-2000202,-2000194,-2000186,-2000178,-2000170,-2000162,-2000154,-2000146,-2000138,-2000130,-2000122,-2000115,-2000107,-2000099,-2000091,-2000083,-2000075,-2000067,-2000059,-2000051,-2000043,-2000035,-2000027,-2000019,-2000011,-2000003,-1999995,-1999987,-1999979,-1999971,-1999963,-1999955,-1999947,-1999939,-1999931,-1999923,-1999915,-1999907,-1999899,-1999891,-1999884,-1999876,-1999868,-1999860,-1999852,-1999844,-1999836,-1999828,-1999820,-1999812,-1999804,-1999796,-1999788,-1999780,-1999772,-1999764,-1999756,-1999748,-1999740,-1999732,-1999724,-1999716,-1999708,-1999700,-1999692,-1999684,-1999676,-1999668,-1999660,-1999652,-1999644,-1999636,-1999628,-1999620,-1999612,-1999604,-1999596,-1999588,-1999580,-1999572,-1999564,-1999556,-1999548,-1999540,-1999532,-1999524,-1999516,-1999509,-1999501,-1999493,-1999485,-1999477,-1999469,-1999461,-1999453,-1999445,-1999437,-1999429,-1999421,-1999413,-1999405,-1999397,-1999389,-1999381,-1999373,-1999365,-1999357,-1999349,-1999341,-1999333,-1999325,-1999317,-1999309,-1999301,-1999293,-1999285,-1999277,-1999269,-1999261,-1999253,-1999245,-1999237,-1999229,-1999221,-1999213,-1999205,-1999197,-1999189,-1999181,-1999173,-1999165,-1999157,-1999149,-1999141,-1999133,-1999125,-1999117,-1999109,-1999101,-1999093,-1999085,-1999077,-1999069,-1999061,-1999053,-1999045,-1999037,-1999029,-1999021,-1999013,-1999005,-1998997,-1998989,-1998980,-1998972,-1998964,-1998956,-1998948,-1998940,-1998932,-1998924,-1998916,-1998908,-1998900,-1998892,-1998884,-1998876,-1998868,-1998860,-1998852,-1998844,-1998836,-1998828,-1998820,-1998812,-1998804,-1998796,-1998788,-1998780,-1998772,-1998764,-1998756,-1998748,-1998740,-1998732,-1998724,-1998716,-1998708,-1998700,-1998692,-1998684,-1998676,-1998668,-1998660,-1998652,-1998644,-1998636,-1998628,-1998620,-1998612,-1998603,-1998595,-1998587,-1998579,-1998571,-1998563,-1998555,-1998547,-1998539,-1998531,-1998523,-1998515,-1998507,-1998499,-1998491,-1998483,-1998475,-1998467,-1998459,-1998451,-1998443,-1998435,-1998427,-1998419,-1998411,-1998403,-1998395,-1998387,-1998379,-1998370,-1998362,-1998354,-1998346,-1998338,-1998330,-1998322,-1998314,-1998306,-1998298,-1998290,-1998282,-1998274,-1998266,-1998258,-1998250,-1998242,-1998234,-1998226,-1998218,-1998210,-1998202,-1998193,-1998185,-1998177,-1998169,-1998161,-1998153,-1998145,-1998137,-1998129,-1998121,-1998113,-1998105,-1998097,-1998089,-1998081,-1998073,-1998065,-1998057,-1998049,-1998040,-1998032,-1998024,-1998016,-1998008,-1998000,-1997992,-1997984,-1997976,-1997968,-1997960,-1997952,-1997944,-1997936,-1997928,-1997920,-1997912,-1997903,-1997895,-1997887,-1997879,-1997871,-1997863,-1997855,-1997847,-1997839,-1997831,-1997823,-1997815,-1997807,-1997799,-1997791,-1997783,-1997774,-1997766,-1997758,-1997750,-1997742,-1997734,-1997726,-1997718,-1997710,-1997702,-1997694,-1997686,-1997678,-1997670,-1997661,-1997653,-1997645,-1997637,-1997629,-1997621,-1997613,-1997605,-1997597,-1997589,-1997581,-1997573,-1997565,-1997556,-1997548,-1997540,-1997532,-1997524,-1997516,-1997508,-1997500,-1997492,-1997484,-1997476,-1997468,-1997460,-1997451,-1997443,-1997435,-1997427,-1997419,-1997411,-1997403,-1997395,-1997387,-1997379,-1997371,-1997362,-1997354,-1997346,-1997338,-1997330,-1997322,-1997314,-1997306,-1997298,-1997290,-1997282,-1997274,-1997265,-1997257,-1997249,-1997241,-1997233,-1997225,-1997217,-1997209,-1997201,-1997193,-1997184,-1997176,-1997168,-1997160,-1997152,-1997144,-1997136,-1997128,-1997120,-1997112,-1997104,-1997095,-1997087,-1997079,-1997071,-1997063,-1997055,-1997047,-1997039,-1997031,-1997023,-1997014,-1997006,-1996998,-1996990,-1996982,-1996974,-1996966,-1996958,-1996950,-1996941,-1996933,-1996925,-1996917,-1996909,-1996901,-1996893,-1996885,-1996877,-1996868,-1996860,-1996852,-1996844,-1996836,-1996828,-1996820,-1996812,-1996804,-1996795,-1996787,-1996779,-1996771,-1996763,-1996755,-1996747,-1996739,-1996731,-1996722,-1996714,-1996706,-1996698,-1996690,-1996682,-1996674,-1996666,-1996658,-1996649,-1996641,-1996633,-1996625,-1996617,-1996609,-1996601,-1996593,-1996584,-1996576,-1996568,-1996560,-1996552,-1996544,-1996536,-1996528,-1996519,-1996511,-1996503,-1996495,-1996487,-1996479,-1996471,-1996463,-1996454,-1996446,-1996438,-1996430,-1996422,-1996414,-1996406,-1996397,-1996389,-1996381,-1996373,-1996365,-1996357,-1996349,-1996341,-1996332,-1996324,-1996316,-1996308,-1996300,-1996292,-1996284,-1996275,-1996267,-1996259,-1996251,-1996243,-1996235,-1996227,-1996219,-1996210,-1996202,-1996194,-1996186,-1996178,-1996170,-1996162,-1996153,-1996145,-1996137,-1996129,-1996121,-1996113,-1996105,-1996096,-1996088,-1996080,-1996072,-1996064,-1996056,-1996048,-1996039,-1996031,-1996023,-1996015,-1996007,-1995999,-1995990,-1995982,-1995974,-1995966,-1995958,-1995950,-1995942,-1995933,-1995925,-1995917,-1995909,-1995901,-1995893,-1995884,-1995876,-1995868,-1995860,-1995852,-1995844,-1995836,-1995827,-1995819,-1995811,-1995803,-1995795,-1995787,-1995778,-1995770,-1995762,-1995754,-1995746,-1995738,-1995729,-1995721,-1995713,-1995705,-1995697,-1995689,-1995680,-1995672,-1995664,-1995656,-1995648,-1995640,-1995632,-1995623,-1995615,-1995607,-1995599,-1995591,-1995583,-1995574,-1995566,-1995558,-1995550,-1995542,-1995533,-1995525,-1995517,-1995509,-1995501,-1995493,-1995484,-1995476,-1995468,-1995460,-1995452,-1995444,-1995435,-1995427,-1995419,-1995411,-1995403,-1995395,-1995386,-1995378,-1995370,-1995362,-1995354,-1995345,-1995337,-1995329,-1995321,-1995313,-1995305,-1995296,-1995288,-1995280,-1995272,-1995264,-1995255,-1995247,-1995239,-1995231,-1995223,-1995215,-1995206,-1995198,-1995190,-1995182,-1995174,-1995165,-1995157,-1995149,-1995141,-1995133,-1995124,-1995116,-1995108,-1995100,-1995092,-1995084,-1995075,-1995067,-1995059,-1995051,-1995043,-1995034,-1995026,-1995018,-1995010,-1995002,-1994993,-1994985,-1994977,-1994969,-1994961,-1994952,-1994944,-1994936,-1994928,-1994920,-1994911,-1994903,-1994895,-1994887,-1994879,-1994870,-1994862,-1994854,-1994846,-1994838,-1994829,-1994821,-1994813,-1994805,-1994797,-1994788,-1994780,-1994772,-1994764,-1994756,-1994747,-1994739,-1994731,-1994723,-1994715,-1994706,-1994698,-1994690,-1994682,-1994674,-1994665,-1994657,-1994649,-1994641,-1994632,-1994624,-1994616,-1994608,-1994600,-1994591,-1994583,-1994575,-1994567,-1994559,-1994550,-1994542,-1994534,-1994526,-1994517,-1994509,-1994501,-1994493,-1994485,-1994476,-1994468,-1994460,-1994452,-1994444,-1994435,-1994427,-1994419,-1994411,-1994402,-1994394,-1994386,-1994378,-1994370,-1994361,-1994353,-1994345,-1994337,-1994328,-1994320,-1994312,-1994304,-1994295,-1994287,-1994279,-1994271,-1994263,-1994254,-1994246,-1994238,-1994230,-1994221,-1994213,-1994205,-1994197,-1994189,-1994180,-1994172,-1994164,-1994156,-1994147,-1994139,-1994131,-1994123,-1994114,-1994106,-1994098,-1994090,-1994081,-1994073,-1994065,-1994057,-1994049,-1994040,-1994032,-1994024,-1994016,-1994007,-1993999,-1993991,-1993983,-1993974,-1993966,-1993958,-1993950,-1993941,-1993933,-1993925,-1993917,-1993908,-1993900,-1993892,-1993884,-1993875,-1993867,-1993859,-1993851,-1993842,-1993834,-1993826,-1993818,-1993809,-1993801,-1993793,-1993785,-1993776,-1993768,-1993760,-1993752,-1993743,-1993735,-1993727,-1993719,-1993710,-1993702,-1993694,-1993686,-1993677,-1993669,-1993661,-1993653,-1993644,-1993636,-1993628,-1993620,-1993611,-1993603,-1993595,-1993587,-1993578,-1993570,-1993562,-1993554,-1993545,-1993537,-1993529,-1993521,-1993512,-1993504,-1993496,-1993488,-1993479,-1993471,-1993463,-1993454,-1993446,-1993438,-1993430,-1993421,-1993413,-1993405,-1993397,-1993388,-1993380,-1993372,-1993364,-1993355,-1993347,-1993339,-1993330,-1993322,-1993314,-1993306,-1993297,-1993289,-1993281,-1993273,-1993264,-1993256,-1993248,-1993239,-1993231,-1993223,-1993215,-1993206,-1993198,-1993190,-1993182,-1993173,-1993165,-1993157,-1993148,-1993140,-1993132,-1993124,-1993115,-1993107,-1993099,-1993090,-1993082,-1993074,-1993066,-1993057,-1993049,-1993041,-1993032,-1993024,-1993016,-1993008,-1992999,-1992991,-1992983,-1992974,-1992966,-1992958,-1992950,-1992941,-1992933,-1992925,-1992916,-1992908,-1992900,-1992892,-1992883,-1992875,-1992867,-1992858,-1992850,-1992842,-1992834,-1992825,-1992817,-1992809,-1992800,-1992792,-1992784,-1992776,-1992767,-1992759,-1992751,-1992742,-1992734,-1992726,-1992717,-1992709,-1992701,-1992693,-1992684,-1992676,-1992668,-1992659,-1992651,-1992643,-1992634,-1992626,-1992618,-1992610,-1992601,-1992593,-1992585,-1992576,-1992568,-1992560,-1992551,-1992543,-1992535,-1992527,-1992518,-1992510,-1992502,-1992493,-1992485,-1992477,-1992468,-1992460,-1992452,-1992443,-1992435,-1992427,-1992418,-1992410,-1992402,-1992394,-1992385,-1992377,-1992369,-1992360,-1992352,-1992344,-1992335,-1992327,-1992319,-1992310,-1992302,-1992294,-1992285,-1992277,-1992269,-1992261,-1992252,-1992244,-1992236,-1992227,-1992219,-1992211,-1992202,-1992194,-1992186,-1992177,-1992169,-1992161,-1992152,-1992144,-1992136,-1992127,-1992119,-1992111,-1992102,-1992094,-1992086,-1992077,-1992069,-1992061,-1992052,-1992044,-1992036,-1992027,-1992019,-1992011,-1992002,-1991994,-1991986,-1991978,-1991969,-1991961,-1991953,-1991944,-1991936,-1991928,-1991919,-1991911,-1991903,-1991894,-1991886,-1991878,-1991869,-1991861,-1991853,-1991844,-1991836,-1991827,-1991819,-1991811,-1991802,-1991794,-1991786,-1991777,-1991769,-1991761,-1991752,-1991744,-1991736,-1991727,-1991719,-1991711,-1991702,-1991694,-1991686,-1991677,-1991669,-1991661,-1991652,-1991644,-1991636,-1991627,-1991619,-1991611,-1991602,-1991594,-1991586,-1991577,-1991569,-1991561,-1991552,-1991544,-1991535,-1991527,-1991519,-1991510,-1991502,-1991494,-1991485,-1991477,-1991469,-1991460,-1991452,-1991444,-1991435,-1991427,-1991419,-1991410,-1991402,-1991393,-1991385,-1991377,-1991368,-1991360,-1991352,-1991343,-1991335,-1991327,-1991318,-1991310,-1991302,-1991293,-1991285,-1991276,-1991268,-1991260,-1991251,-1991243,-1991235,-1991226,-1991218,-1991210,-1991201,-1991193,-1991184,-1991176,-1991168,-1991159,-1991151,-1991143,-1991134,-1991126,-1991118,-1991109,-1991101,-1991092,-1991084,-1991076,-1991067,-1991059,-1991051,-1991042,-1991034,-1991025,-1991017,-1991009,-1991000,-1990992,-1990984,-1990975,-1990967,-1990958,-1990950,-1990942,-1990933,-1990925,-1990917,-1990908,-1990900,-1990891,-1990883,-1990875,-1990866,-1990858,-1990850,-1990841,-1990833,-1990824,-1990816,-1990808,-1990799,-1990791,-1990782,-1990774,-1990766,-1990757,-1990749,-1990741,-1990732,-1990724,-1990715,-1990707,-1990699,-1990690,-1990682,-1990673,-1990665,-1990657,-1990648,-1990640,-1990632,-1990623,-1990615,-1990606,-1990598,-1990590,-1990581,-1990573,-1990564,-1990556,-1990548,-1990539,-1990531,-1990522,-1990514,-1990506,-1990497,-1990489,-1990480,-1990472,-1990464,-1990455,-1990447,-1990438,-1990430,-1990422,-1990413,-1990405,-1990396,-1990388,-1990380,-1990371,-1990363,-1990354,-1990346,-1990338,-1990329,-1990321,-1990312,-1990304,-1990296,-1990287,-1990279,-1990270,-1990262,-1990254,-1990245,-1990237,-1990228,-1990220,-1990212,-1990203,-1990195,-1990186,-1990178,-1990170,-1990161,-1990153,-1990144,-1990136,-1990127,-1990119,-1990111,-1990102,-1990094,-1990085,-1990077,-1990069,-1990060,-1990052,-1990043,-1990035,-1990026,-1990018,-1990010,-1990001,-1989993,-1989984,-1989976,-1989968,-1989959,-1989951,-1989942,-1989934,-1989925,-1989917,-1989909,-1989900,-1989892,-1989883,-1989875,-1989866,-1989858,-1989850,-1989841,-1989833,-1989824,-1989816,-1989808,-1989799,-1989791,-1989782,-1989774,-1989765,-1989757,-1989749,-1989740,-1989732,-1989723,-1989715,-1989706,-1989698,-1989690,-1989681,-1989673,-1989664,-1989656,-1989647,-1989639,-1989630,-1989622,-1989614,-1989605,-1989597,-1989588,-1989580,-1989571,-1989563,-1989555,-1989546,-1989538,-1989529,-1989521,-1989512,-1989504,-1989495,-1989487,-1989479,-1989470,-1989462,-1989453,-1989445,-1989436,-1989428,-1989420,-1989411,-1989403,-1989394,-1989386,-1989377,-1989369,-1989360,-1989352,-1989344,-1989335,-1989327,-1989318,-1989310,-1989301,-1989293,-1989284,-1989276,-1989267,-1989259,-1989251,-1989242,-1989234,-1989225,-1989217,-1989208,-1989200,-1989191,-1989183,-1989175,-1989166,-1989158,-1989149,-1989141,-1989132,-1989124,-1989115,-1989107,-1989098,-1989090,-1989081,-1989073,-1989065,-1989056,-1989048,-1989039,-1989031,-1989022,-1989014,-1989005,-1988997,-1988988,-1988980,-1988972,-1988963,-1988955,-1988946,-1988938,-1988929,-1988921,-1988912,-1988904,-1988895,-1988887,-1988878,-1988870,-1988861,-1988853,-1988845,-1988836,-1988828,-1988819,-1988811,-1988802,-1988794,-1988785,-1988777,-1988768,-1988760,-1988751,-1988743,-1988734,-1988726,-1988717,-1988709,-1988701,-1988692,-1988684,-1988675,-1988667,-1988658,-1988650,-1988641,-1988633,-1988624,-1988616,-1988607,-1988599,-1988590,-1988582,-1988573,-1988565,-1988556,-1988548,-1988539,-1988531,-1988522,-1988514,-1988505,-1988497,-1988489,-1988480,-1988472,-1988463,-1988455,-1988446,-1988438,-1988429,-1988421,-1988412,-1988404,-1988395,-1988387,-1988378,-1988370,-1988361,-1988353,-1988344,-1988336,-1988327,-1988319,-1988310,-1988302,-1988293,-1988285,-1988276,-1988268,-1988259,-1988251,-1988242,-1988234,-1988225,-1988217,-1988208,-1988200,-1988191,-1988183,-1988174,-1988166,-1988157,-1988149,-1988140,-1988132,-1988123,-1988115,-1988106,-1988098,-1988089,-1988081,-1988072,-1988064,-1988055,-1988047,-1988038,-1988030,-1988021,-1988013,-1988004,-1987996,-1987987,-1987979,-1987970,-1987962,-1987953,-1987945,-1987936,-1987928,-1987919,-1987911,-1987902,-1987894,-1987885,-1987877,-1987868,-1987860,-1987851,-1987843,-1987834,-1987826,-1987817,-1987809,-1987800,-1987792,-1987783,-1987775,-1987766,-1987758,-1987749,-1987740,-1987732,-1987723,-1987715,-1987706,-1987698,-1987689,-1987681,-1987672,-1987664,-1987655,-1987647,-1987638,-1987630,-1987621,-1987613,-1987604,-1987596,-1987587,-1987579,-1987570,-1987562,-1987553,-1987545,-1987536,-1987527,-1987519,-1987510,-1987502,-1987493,-1987485,-1987476,-1987468,-1987459,-1987451,-1987442,-1987434,-1987425,-1987417,-1987408,-1987400,-1987391,-1987382,-1987374,-1987365,-1987357,-1987348,-1987340,-1987331,-1987323,-1987314,-1987306,-1987297,-1987289,-1987280,-1987272,-1987263,-1987254,-1987246,-1987237,-1987229,-1987220,-1987212,-1987203,-1987195,-1987186,-1987178,-1987169,-1987161,-1987152,-1987143,-1987135,-1987126,-1987118,-1987109,-1987101,-1987092,-1987084,-1987075,-1987067,-1987058,-1987049,-1987041,-1987032,-1987024,-1987015,-1987007,-1986998,-1986990,-1986981,-1986973,-1986964,-1986955,-1986947,-1986938,-1986930,-1986921,-1986913,-1986904,-1986896,-1986887,-1986878,-1986870,-1986861,-1986853,-1986844,-1986836,-1986827,-1986819,-1986810,-1986801,-1986793,-1986784,-1986776,-1986767,-1986759,-1986750,-1986742,-1986733,-1986724,-1986716,-1986707,-1986699,-1986690,-1986682,-1986673,-1986664,-1986656,-1986647,-1986639,-1986630,-1986622,-1986613,-1986605,-1986596,-1986587,-1986579,-1986570,-1986562,-1986553,-1986545,-1986536,-1986527,-1986519,-1986510,-1986502,-1986493,-1986485,-1986476,-1986467,-1986459,-1986450,-1986442,-1986433,-1986425,-1986416,-1986407,-1986399,-1986390,-1986382,-1986373,-1986365,-1986356,-1986347,-1986339,-1986330,-1986322,-1986313,-1986305,-1986296,-1986287,-1986279,-1986270,-1986262,-1986253,-1986244,-1986236,-1986227,-1986219,-1986210,-1986202,-1986193,-1986184,-1986176,-1986167,-1986159,-1986150,-1986141,-1986133,-1986124,-1986116,-1986107,-1986099,-1986090,-1986081,-1986073,-1986064,-1986056,-1986047,-1986038,-1986030,-1986021,-1986013,-1986004,-1985995,-1985987,-1985978,-1985970,-1985961,-1985952,-1985944,-1985935,-1985927,-1985918,-1985910,-1985901,-1985892,-1985884,-1985875,-1985867,-1985858,-1985849,-1985841,-1985832,-1985824,-1985815,-1985806,-1985798,-1985789,-1985781,-1985772,-1985763,-1985755,-1985746,-1985738,-1985729,-1985720,-1985712,-1985703,-1985695,-1985686,-1985677,-1985669,-1985660,-1985651,-1985643,-1985634,-1985626,-1985617,-1985608,-1985600,-1985591,-1985583,-1985574,-1985565,-1985557,-1985548,-1985540,-1985531,-1985522,-1985514,-1985505,-1985496,-1985488,-1985479,-1985471,-1985462,-1985453,-1985445,-1985436,-1985428,-1985419,-1985410,-1985402,-1985393,-1985384,-1985376,-1985367,-1985359,-1985350,-1985341,-1985333,-1985324,-1985316,-1985307,-1985298,-1985290,-1985281,-1985272,-1985264,-1985255,-1985247,-1985238,-1985229,-1985221,-1985212,-1985203,-1985195,-1985186,-1985178,-1985169,-1985160,-1985152,-1985143,-1985134,-1985126,-1985117,-1985109,-1985100,-1985091,-1985083,-1985074,-1985065,-1985057,-1985048,-1985039,-1985031,-1985022,-1985014,-1985005,-1984996,-1984988,-1984979,-1984970,-1984962,-1984953,-1984944,-1984936,-1984927,-1984919,-1984910,-1984901,-1984893,-1984884,-1984875,-1984867,-1984858,-1984849,-1984841,-1984832,-1984824,-1984815,-1984806,-1984798,-1984789,-1984780,-1984772,-1984763,-1984754,-1984746,-1984737,-1984728,-1984720,-1984711,-1984703,-1984694,-1984685,-1984677,-1984668,-1984659,-1984651,-1984642,-1984633,-1984625,-1984616,-1984607,-1984599,-1984590,-1984581,-1984573,-1984564,-1984555,-1984547,-1984538,-1984529,-1984521,-1984512,-1984504,-1984495,-1984486,-1984478,-1984469,-1984460,-1984452,-1984443,-1984434,-1984426,-1984417,-1984408,-1984400,-1984391,-1984382,-1984374,-1984365,-1984356,-1984348,-1984339,-1984330,-1984322,-1984313,-1984304,-1984296,-1984287,-1984278,-1984270,-1984261,-1984252,-1984244,-1984235,-1984226,-1984218,-1984209,-1984200,-1984192,-1984183,-1984174,-1984166,-1984157,-1984148,-1984140,-1984131,-1984122,-1984114,-1984105,-1984096,-1984088,-1984079,-1984070,-1984062,-1984053,-1984044,-1984036,-1984027,-1984018,-1984010,-1984001,-1983992,-1983984,-1983975,-1983966,-1983957,-1983949,-1983940,-1983931,-1983923,-1983914,-1983905,-1983897,-1983888,-1983879,-1983871,-1983862,-1983853,-1983845,-1983836,-1983827,-1983819,-1983810,-1983801,-1983793,-1983784,-1983775,-1983766,-1983758,-1983749,-1983740,-1983732,-1983723,-1983714,-1983706,-1983697,-1983688,-1983680,-1983671,-1983662,-1983654,-1983645,-1983636,-1983627,-1983619,-1983610,-1983601,-1983593,-1983584,-1983575,-1983567,-1983558,-1983549,-1983540,-1983532,-1983523,-1983514,-1983506,-1983497,-1983488,-1983480,-1983471,-1983462,-1983453,-1983445,-1983436,-1983427,-1983419,-1983410,-1983401,-1983393,-1983384,-1983375,-1983366,-1983358,-1983349,-1983340,-1983332,-1983323,-1983314,-1983306,-1983297,-1983288,-1983279,-1983271,-1983262,-1983253,-1983245,-1983236,-1983227,-1983218,-1983210,-1983201,-1983192,-1983184,-1983175,-1983166,-1983157,-1983149,-1983140,-1983131,-1983123,-1983114,-1983105,-1983096,-1983088,-1983079,-1983070,-1983062,-1983053,-1983044,-1983035,-1983027,-1983018,-1983009,-1983001,-1982992,-1982983,-1982974,-1982966,-1982957,-1982948,-1982940,-1982931,-1982922,-1982913,-1982905,-1982896,-1982887,-1982878,-1982870,-1982861,-1982852,-1982844,-1982835,-1982826,-1982817,-1982809,-1982800,-1982791,-1982782,-1982774,-1982765,-1982756,-1982748,-1982739,-1982730,-1982721,-1982713,-1982704,-1982695,-1982686,-1982678,-1982669,-1982660,-1982652,-1982643,-1982634,-1982625,-1982617,-1982608,-1982599,-1982590,-1982582,-1982573,-1982564,-1982555,-1982547,-1982538,-1982529,-1982520,-1982512,-1982503,-1982494,-1982485,-1982477,-1982468,-1982459,-1982451,-1982442,-1982433,-1982424,-1982416,-1982407,-1982398,-1982389,-1982381,-1982372,-1982363,-1982354,-1982346,-1982337,-1982328,-1982319,-1982311,-1982302,-1982293,-1982284,-1982276,-1982267,-1982258,-1982249,-1982241,-1982232,-1982223,-1982214,-1982206,-1982197,-1982188,-1982179,-1982171,-1982162,-1982153,-1982144,-1982136,-1982127,-1982118,-1982109,-1982101,-1982092,-1982083,-1982074,-1982065,-1982057,-1982048,-1982039,-1982030,-1982022,-1982013,-1982004,-1981995,-1981987,-1981978,-1981969,-1981960,-1981952,-1981943,-1981934,-1981925,-1981917,-1981908,-1981899,-1981890,-1981881,-1981873,-1981864,-1981855,-1981846,-1981838,-1981829,-1981820,-1981811,-1981803,-1981794,-1981785,-1981776,-1981767,-1981759,-1981750,-1981741,-1981732,-1981724,-1981715,-1981706,-1981697,-1981689,-1981680,-1981671,-1981662,-1981653,-1981645,-1981636,-1981627,-1981618,-1981610,-1981601,-1981592,-1981583,-1981574,-1981566,-1981557,-1981548,-1981539,-1981530,-1981522,-1981513,-1981504,-1981495,-1981487,-1981478,-1981469,-1981460,-1981451,-1981443,-1981434,-1981425,-1981416,-1981408,-1981399,-1981390,-1981381,-1981372,-1981364,-1981355,-1981346,-1981337,-1981328,-1981320,-1981311,-1981302,-1981293,-1981284,-1981276,-1981267,-1981258,-1981249,-1981241,-1981232,-1981223,-1981214,-1981205,-1981197,-1981188,-1981179,-1981170,-1981161,-1981153,-1981144,-1981135,-1981126,-1981117,-1981109,-1981100,-1981091,-1981082,-1981073,-1981065,-1981056,-1981047,-1981038,-1981029,-1981021,-1981012,-1981003,-1980994,-1980985,-1980977,-1980968,-1980959,-1980950,-1980941,-1980933,-1980924,-1980915,-1980906,-1980897,-1980888,-1980880,-1980871,-1980862,-1980853,-1980844,-1980836,-1980827,-1980818,-1980809,-1980800,-1980792,-1980783,-1980774,-1980765,-1980756,-1980747,-1980739,-1980730,-1980721,-1980712,-1980703,-1980695,-1980686,-1980677,-1980668,-1980659,-1980651,-1980642,-1980633,-1980624,-1980615,-1980606,-1980598,-1980589,-1980580,-1980571,-1980562,-1980553,-1980545,-1980536,-1980527,-1980518,-1980509,-1980501,-1980492,-1980483,-1980474,-1980465,-1980456,-1980448,-1980439,-1980430,-1980421,-1980412,-1980403,-1980395,-1980386,-1980377,-1980368,-1980359,-1980350,-1980342,-1980333,-1980324,-1980315,-1980306,-1980297,-1980289,-1980280,-1980271,-1980262,-1980253,-1980244,-1980236,-1980227,-1980218,-1980209,-1980200,-1980191,-1980183,-1980174,-1980165,-1980156,-1980147,-1980138,-1980130,-1980121,-1980112,-1980103,-1980094,-1980085,-1980077,-1980068,-1980059,-1980050,-1980041,-1980032,-1980023,-1980015,-1980006,-1979997,-1979988,-1979979,-1979970,-1979962,-1979953,-1979944,-1979935,-1979926,-1979917,-1979908,-1979900,-1979891,-1979882,-1979873,-1979864,-1979855,-1979847,-1979838,-1979829,-1979820,-1979811,-1979802,-1979793,-1979785,-1979776,-1979767,-1979758,-1979749,-1979740,-1979731,-1979723,-1979714,-1979705,-1979696,-1979687,-1979678,-1979669,-1979661,-1979652,-1979643,-1979634,-1979625,-1979616,-1979607,-1979599,-1979590,-1979581,-1979572,-1979563,-1979554,-1979545,-1979536,-1979528,-1979519,-1979510,-1979501,-1979492,-1979483,-1979474,-1979466,-1979457,-1979448,-1979439,-1979430,-1979421,-1979412,-1979403,-1979395,-1979386,-1979377,-1979368,-1979359,-1979350,-1979341,-1979333,-1979324,-1979315,-1979306,-1979297,-1979288,-1979279,-1979270,-1979262,-1979253,-1979244,-1979235,-1979226,-1979217,-1979208,-1979199,-1979190,-1979182,-1979173,-1979164,-1979155,-1979146,-1979137,-1979128,-1979119,-1979111,-1979102,-1979093,-1979084,-1979075,-1979066,-1979057,-1979048,-1979039,-1979031,-1979022,-1979013,-1979004,-1978995,-1978986,-1978977,-1978968,-1978960,-1978951,-1978942,-1978933,-1978924,-1978915,-1978906,-1978897,-1978888,-1978879,-1978871,-1978862,-1978853,-1978844,-1978835,-1978826,-1978817,-1978808,-1978799,-1978791,-1978782,-1978773,-1978764,-1978755,-1978746,-1978737,-1978728,-1978719,-1978710,-1978702,-1978693,-1978684,-1978675,-1978666,-1978657,-1978648,-1978639,-1978630,-1978621,-1978613,-1978604,-1978595,-1978586,-1978577,-1978568,-1978559,-1978550,-1978541,-1978532,-1978524,-1978515,-1978506,-1978497,-1978488,-1978479,-1978470,-1978461,-1978452,-1978443,-1978434,-1978426,-1978417,-1978408,-1978399,-1978390,-1978381,-1978372,-1978363,-1978354,-1978345,-1978336,-1978327,-1978319,-1978310,-1978301,-1978292,-1978283,-1978274,-1978265,-1978256,-1978247,-1978238,-1978229,-1978220,-1978212,-1978203,-1978194,-1978185,-1978176,-1978167,-1978158,-1978149,-1978140,-1978131,-1978122,-1978113,-1978105,-1978096,-1978087,-1978078,-1978069,-1978060,-1978051,-1978042,-1978033,-1978024,-1978015,-1978006,-1977997,-1977988,-1977980,-1977971,-1977962,-1977953,-1977944,-1977935,-1977926,-1977917,-1977908,-1977899,-1977890,-1977881,-1977872,-1977863,-1977854,-1977846,-1977837,-1977828,-1977819,-1977810,-1977801,-1977792,-1977783,-1977774,-1977765,-1977756,-1977747,-1977738,-1977729,-1977720,-1977712,-1977703,-1977694,-1977685,-1977676,-1977667,-1977658,-1977649,-1977640,-1977631,-1977622,-1977613,-1977604,-1977595,-1977586,-1977577,-1977568,-1977559,-1977551,-1977542,-1977533,-1977524,-1977515,-1977506,-1977497,-1977488,-1977479,-1977470,-1977461,-1977452,-1977443,-1977434,-1977425,-1977416,-1977407,-1977398,-1977389,-1977380,-1977372,-1977363,-1977354,-1977345,-1977336,-1977327,-1977318,-1977309,-1977300,-1977291,-1977282,-1977273,-1977264,-1977255,-1977246,-1977237,-1977228,-1977219,-1977210,-1977201,-1977192,-1977183,-1977174,-1977165,-1977157,-1977148,-1977139,-1977130,-1977121,-1977112,-1977103,-1977094,-1977085,-1977076,-1977067,-1977058,-1977049,-1977040,-1977031,-1977022,-1977013,-1977004,-1976995,-1976986,-1976977,-1976968,-1976959,-1976950,-1976941,-1976932,-1976923,-1976914,-1976905,-1976896,-1976887,-1976878,-1976870,-1976861,-1976852,-1976843,-1976834,-1976825,-1976816,-1976807,-1976798,-1976789,-1976780,-1976771,-1976762,-1976753,-1976744,-1976735,-1976726,-1976717,-1976708,-1976699,-1976690,-1976681,-1976672,-1976663,-1976654,-1976645,-1976636,-1976627,-1976618,-1976609,-1976600,-1976591,-1976582,-1976573,-1976564,-1976555,-1976546,-1976537,-1976528,-1976519,-1976510,-1976501,-1976492,-1976483,-1976474,-1976465,-1976456,-1976447,-1976438,-1976429,-1976420,-1976411,-1976402,-1976393,-1976384,-1976375,-1976366,-1976357,-1976348,-1976339,-1976330,-1976321,-1976312,-1976303,-1976294,-1976285,-1976276,-1976267,-1976258,-1976249,-1976240,-1976231,-1976222,-1976213,-1976204,-1976195,-1976186,-1976177,-1976168,-1976159,-1976150,-1976141,-1976132,-1976123,-1976114,-1976105,-1976096,-1976087,-1976078,-1976069,-1976060,-1976051,-1976042,-1976033,-1976024,-1976015,-1976006,-1975997,-1975988,-1975979,-1975970,-1975961,-1975952,-1975943,-1975934,-1975925,-1975916,-1975907,-1975898,-1975889,-1975880,-1975871,-1975862,-1975853,-1975844,-1975835,-1975826,-1975817,-1975808,-1975799,-1975790,-1975781,-1975772,-1975763,-1975754,-1975745,-1975736,-1975727,-1975718,-1975709,-1975700,-1975691,-1975682,-1975673,-1975664,-1975655,-1975646,-1975637,-1975628,-1975618,-1975609,-1975600,-1975591,-1975582,-1975573,-1975564,-1975555,-1975546,-1975537,-1975528,-1975519,-1975510,-1975501,-1975492,-1975483,-1975474,-1975465,-1975456,-1975447,-1975438,-1975429,-1975420,-1975411,-1975402,-1975393,-1975384,-1975375,-1975366,-1975357,-1975348,-1975339,-1975329,-1975320,-1975311,-1975302,-1975293,-1975284,-1975275,-1975266,-1975257,-1975248,-1975239,-1975230,-1975221,-1975212,-1975203,-1975194,-1975185,-1975176,-1975167,-1975158,-1975149,-1975140,-1975131,-1975122,-1975112,-1975103,-1975094,-1975085,-1975076,-1975067,-1975058,-1975049,-1975040,-1975031,-1975022,-1975013,-1975004,-1974995,-1974986,-1974977,-1974968,-1974959,-1974950,-1974941,-1974931,-1974922,-1974913,-1974904,-1974895,-1974886,-1974877,-1974868,-1974859,-1974850,-1974841,-1974832,-1974823,-1974814,-1974805,-1974796,-1974787,-1974778,-1974768,-1974759,-1974750,-1974741,-1974732,-1974723,-1974714,-1974705,-1974696,-1974687,-1974678,-1974669,-1974660,-1974651,-1974642,-1974633,-1974623,-1974614,-1974605,-1974596,-1974587,-1974578,-1974569,-1974560,-1974551,-1974542,-1974533,-1974524,-1974515,-1974506,-1974496,-1974487,-1974478,-1974469,-1974460,-1974451,-1974442,-1974433,-1974424,-1974415,-1974406,-1974397,-1974388,-1974379,-1974369,-1974360,-1974351,-1974342,-1974333,-1974324,-1974315,-1974306,-1974297,-1974288,-1974279,-1974270,-1974261,-1974251,-1974242,-1974233,-1974224,-1974215,-1974206,-1974197,-1974188,-1974179,-1974170,-1974161,-1974152,-1974142,-1974133,-1974124,-1974115,-1974106,-1974097,-1974088,-1974079,-1974070,-1974061,-1974052,-1974042,-1974033,-1974024,-1974015,-1974006,-1973997,-1973988,-1973979,-1973970,-1973961,-1973952,-1973942,-1973933,-1973924,-1973915,-1973906,-1973897,-1973888,-1973879,-1973870,-1973861,-1973852,-1973842,-1973833,-1973824,-1973815,-1973806,-1973797,-1973788,-1973779,-1973770,-1973761,-1973751,-1973742,-1973733,-1973724,-1973715,-1973706,-1973697,-1973688,-1973679,-1973669,-1973660,-1973651,-1973642,-1973633,-1973624,-1973615,-1973606,-1973597,-1973588,-1973578,-1973569,-1973560,-1973551,-1973542,-1973533,-1973524,-1973515,-1973506,-1973496,-1973487,-1973478,-1973469,-1973460,-1973451,-1973442,-1973433,-1973424,-1973414,-1973405,-1973396,-1973387,-1973378,-1973369,-1973360,-1973351,-1973341,-1973332,-1973323,-1973314,-1973305,-1973296,-1973287,-1973278,-1973269,-1973259,-1973250,-1973241,-1973232,-1973223,-1973214,-1973205,-1973196,-1973186,-1973177,-1973168,-1973159,-1973150,-1973141,-1973132,-1973123,-1973113,-1973104,-1973095,-1973086,-1973077,-1973068,-1973059,-1973050,-1973040,-1973031,-1973022,-1973013,-1973004,-1972995,-1972986,-1972976,-1972967,-1972958,-1972949,-1972940,-1972931,-1972922,-1972913,-1972903,-1972894,-1972885,-1972876,-1972867,-1972858,-1972849,-1972839,-1972830,-1972821,-1972812,-1972803,-1972794,-1972785,-1972775,-1972766,-1972757,-1972748,-1972739,-1972730,-1972721,-1972711,-1972702,-1972693,-1972684,-1972675,-1972666,-1972657,-1972647,-1972638,-1972629,-1972620,-1972611,-1972602,-1972593,-1972583,-1972574,-1972565,-1972556,-1972547,-1972538,-1972529,-1972519,-1972510,-1972501,-1972492,-1972483,-1972474,-1972464,-1972455,-1972446,-1972437,-1972428,-1972419,-1972410,-1972400,-1972391,-1972382,-1972373,-1972364,-1972355,-1972345,-1972336,-1972327,-1972318,-1972309,-1972300,-1972291,-1972281,-1972272,-1972263,-1972254,-1972245,-1972236,-1972226,-1972217,-1972208,-1972199,-1972190,-1972181,-1972171,-1972162,-1972153,-1972144,-1972135,-1972126,-1972116,-1972107,-1972098,-1972089,-1972080,-1972071,-1972061,-1972052,-1972043,-1972034,-1972025,-1972016,-1972006,-1971997,-1971988,-1971979,-1971970,-1971961,-1971951,-1971942,-1971933,-1971924,-1971915,-1971905,-1971896,-1971887,-1971878,-1971869,-1971860,-1971850,-1971841,-1971832,-1971823,-1971814,-1971805,-1971795,-1971786,-1971777,-1971768,-1971759,-1971749,-1971740,-1971731,-1971722,-1971713,-1971704,-1971694,-1971685,-1971676,-1971667,-1971658,-1971648,-1971639,-1971630,-1971621,-1971612,-1971602,-1971593,-1971584,-1971575,-1971566,-1971557,-1971547,-1971538,-1971529,-1971520,-1971511,-1971501,-1971492,-1971483,-1971474,-1971465,-1971455,-1971446,-1971437,-1971428,-1971419,-1971409,-1971400,-1971391,-1971382,-1971373,-1971363,-1971354,-1971345,-1971336,-1971327,-1971317,-1971308,-1971299,-1971290,-1971281,-1971271,-1971262,-1971253,-1971244,-1971235,-1971225,-1971216,-1971207,-1971198,-1971189,-1971179,-1971170,-1971161,-1971152,-1971143,-1971133,-1971124,-1971115,-1971106,-1971097,-1971087,-1971078,-1971069,-1971060,-1971051,-1971041,-1971032,-1971023,-1971014,-1971005,-1970995,-1970986,-1970977,-1970968,-1970958,-1970949,-1970940,-1970931,-1970922,-1970912,-1970903,-1970894,-1970885,-1970876,-1970866,-1970857,-1970848,-1970839,-1970829,-1970820,-1970811,-1970802,-1970793,-1970783,-1970774,-1970765,-1970756,-1970746,-1970737,-1970728,-1970719,-1970710,-1970700,-1970691,-1970682,-1970673,-1970663,-1970654,-1970645,-1970636,-1970627,-1970617,-1970608,-1970599,-1970590,-1970580,-1970571,-1970562,-1970553,-1970543,-1970534,-1970525,-1970516,-1970507,-1970497,-1970488,-1970479,-1970470,-1970460,-1970451,-1970442,-1970433,-1970423,-1970414,-1970405,-1970396,-1970387,-1970377,-1970368,-1970359,-1970350,-1970340,-1970331,-1970322,-1970313,-1970303,-1970294,-1970285,-1970276,-1970266,-1970257,-1970248,-1970239,-1970229,-1970220,-1970211,-1970202,-1970192,-1970183,-1970174,-1970165,-1970156,-1970146,-1970137,-1970128,-1970119,-1970109,-1970100,-1970091,-1970082,-1970072,-1970063,-1970054,-1970045,-1970035,-1970026,-1970017,-1970008,-1969998,-1969989,-1969980,-1969971,-1969961,-1969952,-1969943,-1969934,-1969924,-1969915,-1969906,-1969897,-1969887,-1969878,-1969869,-1969859,-1969850,-1969841,-1969832,-1969822,-1969813,-1969804,-1969795,-1969785,-1969776,-1969767,-1969758,-1969748,-1969739,-1969730,-1969721,-1969711,-1969702,-1969693,-1969684,-1969674,-1969665,-1969656,-1969646,-1969637,-1969628,-1969619,-1969609,-1969600,-1969591,-1969582,-1969572,-1969563,-1969554,-1969545,-1969535,-1969526,-1969517,-1969507,-1969498,-1969489,-1969480,-1969470,-1969461,-1969452,-1969443,-1969433,-1969424,-1969415,-1969405,-1969396,-1969387,-1969378,-1969368,-1969359,-1969350,-1969341,-1969331,-1969322,-1969313,-1969303,-1969294,-1969285,-1969276,-1969266,-1969257,-1969248,-1969238,-1969229,-1969220,-1969211,-1969201,-1969192,-1969183,-1969173,-1969164,-1969155,-1969146,-1969136,-1969127,-1969118,-1969108,-1969099,-1969090,-1969081,-1969071,-1969062,-1969053,-1969043,-1969034,-1969025,-1969016,-1969006,-1968997,-1968988,-1968978,-1968969,-1968960,-1968951,-1968941,-1968932,-1968923,-1968913,-1968904,-1968895,-1968886,-1968876,-1968867,-1968858,-1968848,-1968839,-1968830,-1968820,-1968811,-1968802,-1968793,-1968783,-1968774,-1968765,-1968755,-1968746,-1968737,-1968727,-1968718,-1968709,-1968700,-1968690,-1968681,-1968672,-1968662,-1968653,-1968644,-1968634,-1968625,-1968616,-1968606,-1968597,-1968588,-1968579,-1968569,-1968560,-1968551,-1968541,-1968532,-1968523,-1968513,-1968504,-1968495,-1968485,-1968476,-1968467,-1968458,-1968448,-1968439,-1968430,-1968420,-1968411,-1968402,-1968392,-1968383,-1968374,-1968364,-1968355,-1968346,-1968336,-1968327,-1968318,-1968309,-1968299,-1968290,-1968281,-1968271,-1968262,-1968253,-1968243,-1968234,-1968225,-1968215,-1968206,-1968197,-1968187,-1968178,-1968169,-1968159,-1968150,-1968141,-1968131,-1968122,-1968113,-1968103,-1968094,-1968085,-1968075,-1968066,-1968057,-1968047,-1968038,-1968029,-1968019,-1968010,-1968001,-1967991,-1967982,-1967973,-1967963,-1967954,-1967945,-1967935,-1967926,-1967917,-1967907,-1967898,-1967889,-1967879,-1967870,-1967861,-1967851,-1967842,-1967833,-1967823,-1967814,-1967805,-1967795,-1967786,-1967777,-1967767,-1967758,-1967749,-1967739,-1967730,-1967721,-1967711,-1967702,-1967693,-1967683,-1967674,-1967665,-1967655,-1967646,-1967637,-1967627,-1967618,-1967609,-1967599,-1967590,-1967581,-1967571,-1967562,-1967553,-1967543,-1967534,-1967525,-1967515,-1967506,-1967496,-1967487,-1967478,-1967468,-1967459,-1967450,-1967440,-1967431,-1967422,-1967412,-1967403,-1967394,-1967384,-1967375,-1967366,-1967356,-1967347,-1967337,-1967328,-1967319,-1967309,-1967300,-1967291,-1967281,-1967272,-1967263,-1967253,-1967244,-1967235,-1967225,-1967216,-1967206,-1967197,-1967188,-1967178,-1967169,-1967160,-1967150,-1967141,-1967132,-1967122,-1967113,-1967103,-1967094,-1967085,-1967075,-1967066,-1967057,-1967047,-1967038,-1967029,-1967019,-1967010,-1967000,-1966991,-1966982,-1966972,-1966963,-1966954,-1966944,-1966935,-1966925,-1966916,-1966907,-1966897,-1966888,-1966879,-1966869,-1966860,-1966850,-1966841,-1966832,-1966822,-1966813,-1966804,-1966794,-1966785,-1966775,-1966766,-1966757,-1966747,-1966738,-1966729,-1966719,-1966710,-1966700,-1966691,-1966682,-1966672,-1966663,-1966654,-1966644,-1966635,-1966625,-1966616,-1966607,-1966597,-1966588,-1966578,-1966569,-1966560,-1966550,-1966541,-1966531,-1966522,-1966513,-1966503,-1966494,-1966485,-1966475,-1966466,-1966456,-1966447,-1966438,-1966428,-1966419,-1966409,-1966400,-1966391,-1966381,-1966372,-1966362,-1966353,-1966344,-1966334,-1966325,-1966315,-1966306,-1966297,-1966287,-1966278,-1966269,-1966259,-1966250,-1966240,-1966231,-1966222,-1966212,-1966203,-1966193,-1966184,-1966175,-1966165,-1966156,-1966146,-1966137,-1966127,-1966118,-1966109,-1966099,-1966090,-1966080,-1966071,-1966062,-1966052,-1966043,-1966033,-1966024,-1966015,-1966005,-1965996,-1965986,-1965977,-1965968,-1965958,-1965949,-1965939,-1965930,-1965921,-1965911,-1965902,-1965892,-1965883,-1965873,-1965864,-1965855,-1965845,-1965836,-1965826,-1965817,-1965808,-1965798,-1965789,-1965779,-1965770,-1965760,-1965751,-1965742,-1965732,-1965723,-1965713,-1965704,-1965695,-1965685,-1965676,-1965666,-1965657,-1965647,-1965638,-1965629,-1965619,-1965610,-1965600,-1965591,-1965582,-1965572,-1965563,-1965553,-1965544,-1965534,-1965525,-1965516,-1965506,-1965497,-1965487,-1965478,-1965468,-1965459,-1965450,-1965440,-1965431,-1965421,-1965412,-1965402,-1965393,-1965384,-1965374,-1965365,-1965355,-1965346,-1965336,-1965327,-1965317,-1965308,-1965299,-1965289,-1965280,-1965270,-1965261,-1965251,-1965242,-1965233,-1965223,-1965214,-1965204,-1965195,-1965185,-1965176,-1965166,-1965157,-1965148,-1965138,-1965129,-1965119,-1965110,-1965100,-1965091,-1965082,-1965072,-1965063,-1965053,-1965044,-1965034,-1965025,-1965015,-1965006,-1964996,-1964987,-1964978,-1964968,-1964959,-1964949,-1964940,-1964930,-1964921,-1964911,-1964902,-1964893,-1964883,-1964874,-1964864,-1964855,-1964845,-1964836,-1964826,-1964817,-1964807,-1964798,-1964789,-1964779,-1964770,-1964760,-1964751,-1964741,-1964732,-1964722,-1964713,-1964703,-1964694,-1964685,-1964675,-1964666,-1964656,-1964647,-1964637,-1964628,-1964618,-1964609,-1964599,-1964590,-1964580,-1964571,-1964562,-1964552,-1964543,-1964533,-1964524,-1964514,-1964505,-1964495,-1964486,-1964476,-1964467,-1964457,-1964448,-1964438,-1964429,-1964420,-1964410,-1964401,-1964391,-1964382,-1964372,-1964363,-1964353,-1964344,-1964334,-1964325,-1964315,-1964306,-1964296,-1964287,-1964277,-1964268,-1964259,-1964249,-1964240,-1964230,-1964221,-1964211,-1964202,-1964192,-1964183,-1964173,-1964164,-1964154,-1964145,-1964135,-1964126,-1964116,-1964107,-1964097,-1964088,-1964078,-1964069,-1964059,-1964050,-1964040,-1964031,-1964022,-1964012,-1964003,-1963993,-1963984,-1963974,-1963965,-1963955,-1963946,-1963936,-1963927,-1963917,-1963908,-1963898,-1963889,-1963879,-1963870,-1963860,-1963851,-1963841,-1963832,-1963822,-1963813,-1963803,-1963794,-1963784,-1963775,-1963765,-1963756,-1963746,-1963737,-1963727,-1963718,-1963708,-1963699,-1963689,-1963680,-1963670,-1963661,-1963651,-1963642,-1963632,-1963623,-1963613,-1963604,-1963594,-1963585,-1963575,-1963566,-1963556,-1963547,-1963537,-1963528,-1963518,-1963509,-1963499,-1963490,-1963480,-1963471,-1963461,-1963452,-1963442,-1963433,-1963423,-1963414,-1963404,-1963395,-1963385,-1963376,-1963366,-1963357,-1963347,-1963338,-1963328,-1963319,-1963309,-1963300,-1963290,-1963281,-1963271,-1963262,-1963252,-1963243,-1963233,-1963224,-1963214,-1963204,-1963195,-1963185,-1963176,-1963166,-1963157,-1963147,-1963138,-1963128,-1963119,-1963109,-1963100,-1963090,-1963081,-1963071,-1963062,-1963052,-1963043,-1963033,-1963024,-1963014,-1963005,-1962995,-1962986,-1962976,-1962966,-1962957,-1962947,-1962938,-1962928,-1962919,-1962909,-1962900,-1962890,-1962881,-1962871,-1962862,-1962852,-1962843,-1962833,-1962824,-1962814,-1962804,-1962795,-1962785,-1962776,-1962766,-1962757,-1962747,-1962738,-1962728,-1962719,-1962709,-1962700,-1962690,-1962681,-1962671,-1962661,-1962652,-1962642,-1962633,-1962623,-1962614,-1962604,-1962595,-1962585,-1962576,-1962566,-1962557,-1962547,-1962537,-1962528,-1962518,-1962509,-1962499,-1962490,-1962480,-1962471,-1962461,-1962452,-1962442,-1962432,-1962423,-1962413,-1962404,-1962394,-1962385,-1962375,-1962366,-1962356,-1962347,-1962337,-1962327,-1962318,-1962308,-1962299,-1962289,-1962280,-1962270,-1962261,-1962251,-1962242,-1962232,-1962222,-1962213,-1962203,-1962194,-1962184,-1962175,-1962165,-1962156,-1962146,-1962136,-1962127,-1962117,-1962108,-1962098,-1962089,-1962079,-1962070,-1962060,-1962050,-1962041,-1962031,-1962022,-1962012,-1962003,-1961993,-1961983,-1961974,-1961964,-1961955,-1961945,-1961936,-1961926,-1961917,-1961907,-1961897,-1961888,-1961878,-1961869,-1961859,-1961850,-1961840,-1961830,-1961821,-1961811,-1961802,-1961792,-1961783,-1961773,-1961763,-1961754,-1961744,-1961735,-1961725,-1961716,-1961706,-1961696,-1961687,-1961677,-1961668,-1961658,-1961649,-1961639,-1961629,-1961620,-1961610,-1961601,-1961591,-1961582,-1961572,-1961562,-1961553,-1961543,-1961534,-1961524,-1961514,-1961505,-1961495,-1961486,-1961476,-1961467,-1961457,-1961447,-1961438,-1961428,-1961419,-1961409,-1961399,-1961390,-1961380,-1961371,-1961361,-1961352,-1961342,-1961332,-1961323,-1961313,-1961304,-1961294,-1961284,-1961275,-1961265,-1961256,-1961246,-1961236,-1961227,-1961217,-1961208,-1961198,-1961188,-1961179,-1961169,-1961160,-1961150,-1961141,-1961131,-1961121,-1961112,-1961102,-1961093,-1961083,-1961073,-1961064,-1961054,-1961045,-1961035,-1961025,-1961016,-1961006,-1960997,-1960987,-1960977,-1960968,-1960958,-1960949,-1960939,-1960929,-1960920,-1960910,-1960901,-1960891,-1960881,-1960872,-1960862,-1960853,-1960843,-1960833,-1960824,-1960814,-1960804,-1960795,-1960785,-1960776,-1960766,-1960756,-1960747,-1960737,-1960728,-1960718,-1960708,-1960699,-1960689,-1960680,-1960670,-1960660,-1960651,-1960641,-1960631,-1960622,-1960612,-1960603,-1960593,-1960583,-1960574,-1960564,-1960555,-1960545,-1960535,-1960526,-1960516,-1960506,-1960497,-1960487,-1960478,-1960468,-1960458,-1960449,-1960439,-1960430,-1960420,-1960410,-1960401,-1960391,-1960381,-1960372,-1960362,-1960353,-1960343,-1960333,-1960324,-1960314,-1960304,-1960295,-1960285,-1960276,-1960266,-1960256,-1960247,-1960237,-1960227,-1960218,-1960208,-1960198,-1960189,-1960179,-1960170,-1960160,-1960150,-1960141,-1960131,-1960121,-1960112,-1960102,-1960093,-1960083,-1960073,-1960064,-1960054,-1960044,-1960035,-1960025,-1960015,-1960006,-1959996,-1959987,-1959977,-1959967,-1959958,-1959948,-1959938,-1959929,-1959919,-1959909,-1959900,-1959890,-1959880,-1959871,-1959861,-1959852,-1959842,-1959832,-1959823,-1959813,-1959803,-1959794,-1959784,-1959774,-1959765,-1959755,-1959745,-1959736,-1959726,-1959717,-1959707,-1959697,-1959688,-1959678,-1959668,-1959659,-1959649,-1959639,-1959630,-1959620,-1959610,-1959601,-1959591,-1959581,-1959572,-1959562,-1959552,-1959543,-1959533,-1959523,-1959514,-1959504,-1959494,-1959485,-1959475,-1959466,-1959456,-1959446,-1959437,-1959427,-1959417,-1959408,-1959398,-1959388,-1959379,-1959369,-1959359,-1959350,-1959340,-1959330,-1959321,-1959311,-1959301,-1959292,-1959282,-1959272,-1959263,-1959253,-1959243,-1959234,-1959224,-1959214,-1959205,-1959195,-1959185,-1959176,-1959166,-1959156,-1959147,-1959137,-1959127,-1959118,-1959108,-1959098,-1959089,-1959079,-1959069,-1959060,-1959050,-1959040,-1959031,-1959021,-1959011,-1959002,-1958992,-1958982,-1958972,-1958963,-1958953,-1958943,-1958934,-1958924,-1958914,-1958905,-1958895,-1958885,-1958876,-1958866,-1958856,-1958847,-1958837,-1958827,-1958818,-1958808,-1958798,-1958789,-1958779,-1958769,-1958759,-1958750,-1958740,-1958730,-1958721,-1958711,-1958701,-1958692,-1958682,-1958672,-1958663,-1958653,-1958643,-1958634,-1958624,-1958614,-1958604,-1958595,-1958585,-1958575,-1958566,-1958556,-1958546,-1958537,-1958527,-1958517,-1958508,-1958498,-1958488,-1958478,-1958469,-1958459,-1958449,-1958440,-1958430,-1958420,-1958411,-1958401,-1958391,-1958382,-1958372,-1958362,-1958352,-1958343,-1958333,-1958323,-1958314,-1958304,-1958294,-1958285,-1958275,-1958265,-1958255,-1958246,-1958236,-1958226,-1958217,-1958207,-1958197,-1958187,-1958178,-1958168,-1958158,-1958149,-1958139,-1958129,-1958120,-1958110,-1958100,-1958090,-1958081,-1958071,-1958061,-1958052,-1958042,-1958032,-1958022,-1958013,-1958003,-1957993,-1957984,-1957974,-1957964,-1957954,-1957945,-1957935,-1957925,-1957916,-1957906,-1957896,-1957886,-1957877,-1957867,-1957857,-1957848,-1957838,-1957828,-1957818,-1957809,-1957799,-1957789,-1957779,-1957770,-1957760,-1957750,-1957741,-1957731,-1957721,-1957711,-1957702,-1957692,-1957682,-1957673,-1957663,-1957653,-1957643,-1957634,-1957624,-1957614,-1957604,-1957595,-1957585,-1957575,-1957566,-1957556,-1957546,-1957536,-1957527,-1957517,-1957507,-1957497,-1957488,-1957478,-1957468,-1957458,-1957449,-1957439,-1957429,-1957420,-1957410,-1957400,-1957390,-1957381,-1957371,-1957361,-1957351,-1957342,-1957332,-1957322,-1957312,-1957303,-1957293,-1957283,-1957273,-1957264,-1957254,-1957244,-1957234,-1957225,-1957215,-1957205,-1957196,-1957186,-1957176,-1957166,-1957157,-1957147,-1957137,-1957127,-1957118,-1957108,-1957098,-1957088,-1957079,-1957069,-1957059,-1957049,-1957040,-1957030,-1957020,-1957010,-1957001,-1956991,-1956981,-1956971,-1956962,-1956952,-1956942,-1956932,-1956923,-1956913,-1956903,-1956893,-1956884,-1956874,-1956864,-1956854,-1956845,-1956835,-1956825,-1956815,-1956805,-1956796,-1956786,-1956776,-1956766,-1956757,-1956747,-1956737,-1956727,-1956718,-1956708,-1956698,-1956688,-1956679,-1956669,-1956659,-1956649,-1956640,-1956630,-1956620,-1956610,-1956600,-1956591,-1956581,-1956571,-1956561,-1956552,-1956542,-1956532,-1956522,-1956513,-1956503,-1956493,-1956483,-1956474,-1956464,-1956454,-1956444,-1956434,-1956425,-1956415,-1956405,-1956395,-1956386,-1956376,-1956366,-1956356,-1956346,-1956337,-1956327,-1956317,-1956307,-1956298,-1956288,-1956278,-1956268,-1956258,-1956249,-1956239,-1956229,-1956219,-1956210,-1956200,-1956190,-1956180,-1956170,-1956161,-1956151,-1956141,-1956131,-1956122,-1956112,-1956102,-1956092,-1956082,-1956073,-1956063,-1956053,-1956043,-1956033,-1956024,-1956014,-1956004,-1955994,-1955985,-1955975,-1955965,-1955955,-1955945,-1955936,-1955926,-1955916,-1955906,-1955896,-1955887,-1955877,-1955867,-1955857,-1955847,-1955838,-1955828,-1955818,-1955808,-1955798,-1955789,-1955779,-1955769,-1955759,-1955750,-1955740,-1955730,-1955720,-1955710,-1955701,-1955691,-1955681,-1955671,-1955661,-1955652,-1955642,-1955632,-1955622,-1955612,-1955603,-1955593,-1955583,-1955573,-1955563,-1955553,-1955544,-1955534,-1955524,-1955514,-1955504,-1955495,-1955485,-1955475,-1955465,-1955455,-1955446,-1955436,-1955426,-1955416,-1955406,-1955397,-1955387,-1955377,-1955367,-1955357,-1955348,-1955338,-1955328,-1955318,-1955308,-1955298,-1955289,-1955279,-1955269,-1955259,-1955249,-1955240,-1955230,-1955220,-1955210,-1955200,-1955190,-1955181,-1955171,-1955161,-1955151,-1955141,-1955132,-1955122,-1955112,-1955102,-1955092,-1955082,-1955073,-1955063,-1955053,-1955043,-1955033,-1955024,-1955014,-1955004,-1954994,-1954984,-1954974,-1954965,-1954955,-1954945,-1954935,-1954925,-1954915,-1954906,-1954896,-1954886,-1954876,-1954866,-1954856,-1954847,-1954837,-1954827,-1954817,-1954807,-1954797,-1954788,-1954778,-1954768,-1954758,-1954748,-1954738,-1954729,-1954719,-1954709,-1954699,-1954689,-1954679,-1954670,-1954660,-1954650,-1954640,-1954630,-1954620,-1954611,-1954601,-1954591,-1954581,-1954571,-1954561,-1954552,-1954542,-1954532,-1954522,-1954512,-1954502,-1954492,-1954483,-1954473,-1954463,-1954453,-1954443,-1954433,-1954424,-1954414,-1954404,-1954394,-1954384,-1954374,-1954364,-1954355,-1954345,-1954335,-1954325,-1954315,-1954305,-1954296,-1954286,-1954276,-1954266,-1954256,-1954246,-1954236,-1954227,-1954217,-1954207,-1954197,-1954187,-1954177,-1954167,-1954158,-1954148,-1954138,-1954128,-1954118,-1954108,-1954098,-1954089,-1954079,-1954069,-1954059,-1954049,-1954039,-1954029,-1954020,-1954010,-1954000,-1953990,-1953980,-1953970,-1953960,-1953951,-1953941,-1953931,-1953921,-1953911,-1953901,-1953891,-1953881,-1953872,-1953862,-1953852,-1953842,-1953832,-1953822,-1953812,-1953803,-1953793,-1953783,-1953773,-1953763,-1953753,-1953743,-1953733,-1953724,-1953714,-1953704,-1953694,-1953684,-1953674,-1953664,-1953654,-1953645,-1953635,-1953625,-1953615,-1953605,-1953595,-1953585,-1953575,-1953566,-1953556,-1953546,-1953536,-1953526,-1953516,-1953506,-1953496,-1953487,-1953477,-1953467,-1953457,-1953447,-1953437,-1953427,-1953417,-1953407,-1953398,-1953388,-1953378,-1953368,-1953358,-1953348,-1953338,-1953328,-1953319,-1953309,-1953299,-1953289,-1953279,-1953269,-1953259,-1953249,-1953239,-1953230,-1953220,-1953210,-1953200,-1953190,-1953180,-1953170,-1953160,-1953150,-1953140,-1953131,-1953121,-1953111,-1953101,-1953091,-1953081,-1953071,-1953061,-1953051,-1953042,-1953032,-1953022,-1953012,-1953002,-1952992,-1952982,-1952972,-1952962,-1952952,-1952943,-1952933,-1952923,-1952913,-1952903,-1952893,-1952883,-1952873,-1952863,-1952853,-1952844,-1952834,-1952824,-1952814,-1952804,-1952794,-1952784,-1952774,-1952764,-1952754,-1952744,-1952735,-1952725,-1952715,-1952705,-1952695,-1952685,-1952675,-1952665,-1952655,-1952645,-1952635,-1952626,-1952616,-1952606,-1952596,-1952586,-1952576,-1952566,-1952556,-1952546,-1952536,-1952526,-1952516,-1952507,-1952497,-1952487,-1952477,-1952467,-1952457,-1952447,-1952437,-1952427,-1952417,-1952407,-1952397,-1952388,-1952378,-1952368,-1952358,-1952348,-1952338,-1952328,-1952318,-1952308,-1952298,-1952288,-1952278,-1952268,-1952259,-1952249,-1952239,-1952229,-1952219,-1952209,-1952199,-1952189,-1952179,-1952169,-1952159,-1952149,-1952139,-1952129,-1952120,-1952110,-1952100,-1952090,-1952080,-1952070,-1952060,-1952050,-1952040,-1952030,-1952020,-1952010,-1952000,-1951990,-1951980,-1951971,-1951961,-1951951,-1951941,-1951931,-1951921,-1951911,-1951901,-1951891,-1951881,-1951871,-1951861,-1951851,-1951841,-1951831,-1951821,-1951811,-1951802,-1951792,-1951782,-1951772,-1951762,-1951752,-1951742,-1951732,-1951722,-1951712,-1951702,-1951692,-1951682,-1951672,-1951662,-1951652,-1951642,-1951632,-1951623,-1951613,-1951603,-1951593,-1951583,-1951573,-1951563,-1951553,-1951543,-1951533,-1951523,-1951513,-1951503,-1951493,-1951483,-1951473,-1951463,-1951453,-1951443,-1951433,-1951423,-1951414,-1951404,-1951394,-1951384,-1951374,-1951364,-1951354,-1951344,-1951334,-1951324,-1951314,-1951304,-1951294,-1951284,-1951274,-1951264,-1951254,-1951244,-1951234,-1951224,-1951214,-1951204,-1951194,-1951184,-1951174,-1951164,-1951155,-1951145,-1951135,-1951125,-1951115,-1951105,-1951095,-1951085,-1951075,-1951065,-1951055,-1951045,-1951035,-1951025,-1951015,-1951005,-1950995,-1950985,-1950975,-1950965,-1950955,-1950945,-1950935,-1950925,-1950915,-1950905,-1950895,-1950885,-1950875,-1950865,-1950855,-1950845,-1950835,-1950825,-1950815,-1950805,-1950795,-1950786,-1950776,-1950766,-1950756,-1950746,-1950736,-1950726,-1950716,-1950706,-1950696,-1950686,-1950676,-1950666,-1950656,-1950646,-1950636,-1950626,-1950616,-1950606,-1950596,-1950586,-1950576,-1950566,-1950556,-1950546,-1950536,-1950526,-1950516,-1950506,-1950496,-1950486,-1950476,-1950466,-1950456,-1950446,-1950436,-1950426,-1950416,-1950406,-1950396,-1950386,-1950376,-1950366,-1950356,-1950346,-1950336,-1950326,-1950316,-1950306,-1950296,-1950286,-1950276,-1950266,-1950256,-1950246,-1950236,-1950226,-1950216,-1950206,-1950196,-1950186,-1950176,-1950166,-1950156,-1950146,-1950136,-1950126,-1950116,-1950106,-1950096,-1950086,-1950076,-1950066,-1950056,-1950046,-1950036,-1950026,-1950016,-1950006,-1949996,-1949986,-1949976,-1949966,-1949956,-1949946,-1949936,-1949926,-1949916,-1949906,-1949896,-1949886,-1949876,-1949866,-1949856,-1949846,-1949836,-1949826,-1949816,-1949806,-1949796,-1949786,-1949776,-1949766,-1949756,-1949746,-1949736,-1949726,-1949716,-1949706,-1949696,-1949686,-1949676,-1949666,-1949656,-1949645,-1949635,-1949625,-1949615,-1949605,-1949595,-1949585,-1949575,-1949565,-1949555,-1949545,-1949535,-1949525,-1949515,-1949505,-1949495,-1949485,-1949475,-1949465,-1949455,-1949445,-1949435,-1949425,-1949415,-1949405,-1949395,-1949385,-1949375,-1949365,-1949355,-1949345,-1949335,-1949325,-1949315,-1949305,-1949295,-1949285,-1949274,-1949264,-1949254,-1949244,-1949234,-1949224,-1949214,-1949204,-1949194,-1949184,-1949174,-1949164,-1949154,-1949144,-1949134,-1949124,-1949114,-1949104,-1949094,-1949084,-1949074,-1949064,-1949054,-1949044,-1949034,-1949024,-1949013,-1949003,-1948993,-1948983,-1948973,-1948963,-1948953,-1948943,-1948933,-1948923,-1948913,-1948903,-1948893,-1948883,-1948873,-1948863,-1948853,-1948843,-1948833,-1948823,-1948813,-1948802,-1948792,-1948782,-1948772,-1948762,-1948752,-1948742,-1948732,-1948722,-1948712,-1948702,-1948692,-1948682,-1948672,-1948662,-1948652,-1948642,-1948632,-1948621,-1948611,-1948601,-1948591,-1948581,-1948571,-1948561,-1948551,-1948541,-1948531,-1948521,-1948511,-1948501,-1948491,-1948481,-1948471,-1948461,-1948450,-1948440,-1948430,-1948420,-1948410,-1948400,-1948390,-1948380,-1948370,-1948360,-1948350,-1948340,-1948330,-1948320,-1948310,-1948299,-1948289,-1948279,-1948269,-1948259,-1948249,-1948239,-1948229,-1948219,-1948209,-1948199,-1948189,-1948179,-1948169,-1948158,-1948148,-1948138,-1948128,-1948118,-1948108,-1948098,-1948088,-1948078,-1948068,-1948058,-1948048,-1948038,-1948027,-1948017,-1948007,-1947997,-1947987,-1947977,-1947967,-1947957,-1947947,-1947937,-1947927,-1947917,-1947906,-1947896,-1947886,-1947876,-1947866,-1947856,-1947846,-1947836,-1947826,-1947816,-1947806,-1947796,-1947785,-1947775,-1947765,-1947755,-1947745,-1947735,-1947725,-1947715,-1947705,-1947695,-1947685,-1947674,-1947664,-1947654,-1947644,-1947634,-1947624,-1947614,-1947604,-1947594,-1947584,-1947574,-1947563,-1947553,-1947543,-1947533,-1947523,-1947513,-1947503,-1947493,-1947483,-1947473,-1947462,-1947452,-1947442,-1947432,-1947422,-1947412,-1947402,-1947392,-1947382,-1947372,-1947361,-1947351,-1947341,-1947331,-1947321,-1947311,-1947301,-1947291,-1947281,-1947270,-1947260,-1947250,-1947240,-1947230,-1947220,-1947210,-1947200,-1947190,-1947180,-1947169,-1947159,-1947149,-1947139,-1947129,-1947119,-1947109,-1947099,-1947089,-1947078,-1947068,-1947058,-1947048,-1947038,-1947028,-1947018,-1947008,-1946997,-1946987,-1946977,-1946967,-1946957,-1946947,-1946937,-1946927,-1946917,-1946906,-1946896,-1946886,-1946876,-1946866,-1946856,-1946846,-1946836,-1946825,-1946815,-1946805,-1946795,-1946785,-1946775,-1946765,-1946755,-1946744,-1946734,-1946724,-1946714,-1946704,-1946694,-1946684,-1946674,-1946663,-1946653,-1946643,-1946633,-1946623,-1946613,-1946603,-1946593,-1946582,-1946572,-1946562,-1946552,-1946542,-1946532,-1946522,-1946511,-1946501,-1946491,-1946481,-1946471,-1946461,-1946451,-1946441,-1946430,-1946420,-1946410,-1946400,-1946390,-1946380,-1946370,-1946359,-1946349,-1946339,-1946329,-1946319,-1946309,-1946299,-1946288,-1946278,-1946268,-1946258,-1946248,-1946238,-1946228,-1946217,-1946207,-1946197,-1946187,-1946177,-1946167,-1946157,-1946146,-1946136,-1946126,-1946116,-1946106,-1946096,-1946086,-1946075,-1946065,-1946055,-1946045,-1946035,-1946025,-1946015,-1946004,-1945994,-1945984,-1945974,-1945964,-1945954,-1945943,-1945933,-1945923,-1945913,-1945903,-1945893,-1945883,-1945872,-1945862,-1945852,-1945842,-1945832,-1945822,-1945811,-1945801,-1945791,-1945781,-1945771,-1945761,-1945750,-1945740,-1945730,-1945720,-1945710,-1945700,-1945689,-1945679,-1945669,-1945659,-1945649,-1945639,-1945628,-1945618,-1945608,-1945598,-1945588,-1945578,-1945567,-1945557,-1945547,-1945537,-1945527,-1945517,-1945506,-1945496,-1945486,-1945476,-1945466,-1945456,-1945445,-1945435,-1945425,-1945415,-1945405,-1945395,-1945384,-1945374,-1945364,-1945354,-1945344,-1945334,-1945323,-1945313,-1945303,-1945293,-1945283,-1945272,-1945262,-1945252,-1945242,-1945232,-1945222,-1945211,-1945201,-1945191,-1945181,-1945171,-1945161,-1945150,-1945140,-1945130,-1945120,-1945110,-1945099,-1945089,-1945079,-1945069,-1945059,-1945048,-1945038,-1945028,-1945018,-1945008,-1944998,-1944987,-1944977,-1944967,-1944957,-1944947,-1944936,-1944926,-1944916,-1944906,-1944896,-1944885,-1944875,-1944865,-1944855,-1944845,-1944835,-1944824,-1944814,-1944804,-1944794,-1944784,-1944773,-1944763,-1944753,-1944743,-1944733,-1944722,-1944712,-1944702,-1944692,-1944682,-1944671,-1944661,-1944651,-1944641,-1944631,-1944620,-1944610,-1944600,-1944590,-1944580,-1944569,-1944559,-1944549,-1944539,-1944529,-1944518,-1944508,-1944498,-1944488,-1944478,-1944467,-1944457,-1944447,-1944437,-1944427,-1944416,-1944406,-1944396,-1944386,-1944375,-1944365,-1944355,-1944345,-1944335,-1944324,-1944314,-1944304,-1944294,-1944284,-1944273,-1944263,-1944253,-1944243,-1944232,-1944222,-1944212,-1944202,-1944192,-1944181,-1944171,-1944161,-1944151,-1944141,-1944130,-1944120,-1944110,-1944100,-1944089,-1944079,-1944069,-1944059,-1944049,-1944038,-1944028,-1944018,-1944008,-1943997,-1943987,-1943977,-1943967,-1943957,-1943946,-1943936,-1943926,-1943916,-1943905,-1943895,-1943885,-1943875,-1943865,-1943854,-1943844,-1943834,-1943824,-1943813,-1943803,-1943793,-1943783,-1943772,-1943762,-1943752,-1943742,-1943732,-1943721,-1943711,-1943701,-1943691,-1943680,-1943670,-1943660,-1943650,-1943639,-1943629,-1943619,-1943609,-1943598,-1943588,-1943578,-1943568,-1943558,-1943547,-1943537,-1943527,-1943517,-1943506,-1943496,-1943486,-1943476,-1943465,-1943455,-1943445,-1943435,-1943424,-1943414,-1943404,-1943394,-1943383,-1943373,-1943363,-1943353,-1943342,-1943332,-1943322,-1943312,-1943301,-1943291,-1943281,-1943271,-1943260,-1943250,-1943240,-1943230,-1943219,-1943209,-1943199,-1943189,-1943178,-1943168,-1943158,-1943148,-1943137,-1943127,-1943117,-1943107,-1943096,-1943086,-1943076,-1943066,-1943055,-1943045,-1943035,-1943025,-1943014,-1943004,-1942994,-1942984,-1942973,-1942963,-1942953,-1942943,-1942932,-1942922,-1942912,-1942902,-1942891,-1942881,-1942871,-1942860,-1942850,-1942840,-1942830,-1942819,-1942809,-1942799,-1942789,-1942778,-1942768,-1942758,-1942748,-1942737,-1942727,-1942717,-1942707,-1942696,-1942686,-1942676,-1942665,-1942655,-1942645,-1942635,-1942624,-1942614,-1942604,-1942594,-1942583,-1942573,-1942563,-1942552,-1942542,-1942532,-1942522,-1942511,-1942501,-1942491,-1942481,-1942470,-1942460,-1942450,-1942439,-1942429,-1942419,-1942409,-1942398,-1942388,-1942378,-1942367,-1942357,-1942347,-1942337,-1942326,-1942316,-1942306,-1942295,-1942285,-1942275,-1942265,-1942254,-1942244,-1942234,-1942223,-1942213,-1942203,-1942193,-1942182,-1942172,-1942162,-1942151,-1942141,-1942131,-1942121,-1942110,-1942100,-1942090,-1942079,-1942069,-1942059,-1942049,-1942038,-1942028,-1942018,-1942007,-1941997,-1941987,-1941977,-1941966,-1941956,-1941946,-1941935,-1941925,-1941915,-1941904,-1941894,-1941884,-1941874,-1941863,-1941853,-1941843,-1941832,-1941822,-1941812,-1941801,-1941791,-1941781,-1941771,-1941760,-1941750,-1941740,-1941729,-1941719,-1941709,-1941698,-1941688,-1941678,-1941668,-1941657,-1941647,-1941637,-1941626,-1941616,-1941606,-1941595,-1941585,-1941575,-1941564,-1941554,-1941544,-1941534,-1941523,-1941513,-1941503,-1941492,-1941482,-1941472,-1941461,-1941451,-1941441,-1941430,-1941420,-1941410,-1941400,-1941389,-1941379,-1941369,-1941358,-1941348,-1941338,-1941327,-1941317,-1941307,-1941296,-1941286,-1941276,-1941265,-1941255,-1941245,-1941234,-1941224,-1941214,-1941203,-1941193,-1941183,-1941173,-1941162,-1941152,-1941142,-1941131,-1941121,-1941111,-1941100,-1941090,-1941080,-1941069,-1941059,-1941049,-1941038,-1941028,-1941018,-1941007,-1940997,-1940987,-1940976,-1940966,-1940956,-1940945,-1940935,-1940925,-1940914,-1940904,-1940894,-1940883,-1940873,-1940863,-1940852,-1940842,-1940832,-1940821,-1940811,-1940801,-1940790,-1940780,-1940770,-1940759,-1940749,-1940739,-1940728,-1940718,-1940708,-1940697,-1940687,-1940677,-1940666,-1940656,-1940646,-1940635,-1940625,-1940615,-1940604,-1940594,-1940584,-1940573,-1940563,-1940553,-1940542,-1940532,-1940521,-1940511,-1940501,-1940490,-1940480,-1940470,-1940459,-1940449,-1940439,-1940428,-1940418,-1940408,-1940397,-1940387,-1940377,-1940366,-1940356,-1940346,-1940335,-1940325,-1940315,-1940304,-1940294,-1940283,-1940273,-1940263,-1940252,-1940242,-1940232,-1940221,-1940211,-1940201,-1940190,-1940180,-1940170,-1940159,-1940149,-1940138,-1940128,-1940118,-1940107,-1940097,-1940087,-1940076,-1940066,-1940056,-1940045,-1940035,-1940025,-1940014,-1940004,-1939993,-1939983,-1939973,-1939962,-1939952,-1939942,-1939931,-1939921,-1939911,-1939900,-1939890,-1939879,-1939869,-1939859,-1939848,-1939838,-1939828,-1939817,-1939807,-1939796,-1939786,-1939776,-1939765,-1939755,-1939745,-1939734,-1939724,-1939713,-1939703,-1939693,-1939682,-1939672,-1939662,-1939651,-1939641,-1939631,-1939620,-1939610,-1939599,-1939589,-1939579,-1939568,-1939558,-1939547,-1939537,-1939527,-1939516,-1939506,-1939496,-1939485,-1939475,-1939464,-1939454,-1939444,-1939433,-1939423,-1939413,-1939402,-1939392,-1939381,-1939371,-1939361,-1939350,-1939340,-1939329,-1939319,-1939309,-1939298,-1939288,-1939278,-1939267,-1939257,-1939246,-1939236,-1939226,-1939215,-1939205,-1939194,-1939184,-1939174,-1939163,-1939153,-1939142,-1939132,-1939122,-1939111,-1939101,-1939090,-1939080,-1939070,-1939059,-1939049,-1939038,-1939028,-1939018,-1939007,-1938997,-1938987,-1938976,-1938966,-1938955,-1938945,-1938935,-1938924,-1938914,-1938903,-1938893,-1938883,-1938872,-1938862,-1938851,-1938841,-1938830,-1938820,-1938810,-1938799,-1938789,-1938778,-1938768,-1938758,-1938747,-1938737,-1938726,-1938716,-1938706,-1938695,-1938685,-1938674,-1938664,-1938654,-1938643,-1938633,-1938622,-1938612,-1938602,-1938591,-1938581,-1938570,-1938560,-1938549,-1938539,-1938529,-1938518,-1938508,-1938497,-1938487,-1938477,-1938466,-1938456,-1938445,-1938435,-1938424,-1938414,-1938404,-1938393,-1938383,-1938372,-1938362,-1938352,-1938341,-1938331,-1938320,-1938310,-1938299,-1938289,-1938279,-1938268,-1938258,-1938247,-1938237,-1938226,-1938216,-1938206,-1938195,-1938185,-1938174,-1938164,-1938153,-1938143,-1938133,-1938122,-1938112,-1938101,-1938091,-1938080,-1938070,-1938060,-1938049,-1938039,-1938028,-1938018,-1938007,-1937997,-1937987,-1937976,-1937966,-1937955,-1937945,-1937934,-1937924,-1937914,-1937903,-1937893,-1937882,-1937872,-1937861,-1937851,-1937841,-1937830,-1937820,-1937809,-1937799,-1937788,-1937778,-1937767,-1937757,-1937747,-1937736,-1937726,-1937715,-1937705,-1937694,-1937684,-1937673,-1937663,-1937653,-1937642,-1937632,-1937621,-1937611,-1937600,-1937590,-1937579,-1937569,-1937559,-1937548,-1937538,-1937527,-1937517,-1937506,-1937496,-1937485,-1937475,-1937465,-1937454,-1937444,-1937433,-1937423,-1937412,-1937402,-1937391,-1937381,-1937370,-1937360,-1937350,-1937339,-1937329,-1937318,-1937308,-1937297,-1937287,-1937276,-1937266,-1937255,-1937245,-1937235,-1937224,-1937214,-1937203,-1937193,-1937182,-1937172,-1937161,-1937151,-1937140,-1937130,-1937119,-1937109,-1937099,-1937088,-1937078,-1937067,-1937057,-1937046,-1937036,-1937025,-1937015,-1937004,-1936994,-1936983,-1936973,-1936962,-1936952,-1936942,-1936931,-1936921,-1936910,-1936900,-1936889,-1936879,-1936868,-1936858,-1936847,-1936837,-1936826,-1936816,-1936805,-1936795,-1936784,-1936774,-1936763,-1936753,-1936743,-1936732,-1936722,-1936711,-1936701,-1936690,-1936680,-1936669,-1936659,-1936648,-1936638,-1936627,-1936617,-1936606,-1936596,-1936585,-1936575,-1936564,-1936554,-1936543,-1936533,-1936522,-1936512,-1936502,-1936491,-1936481,-1936470,-1936460,-1936449,-1936439,-1936428,-1936418,-1936407,-1936397,-1936386,-1936376,-1936365,-1936355,-1936344,-1936334,-1936323,-1936313,-1936302,-1936292,-1936281,-1936271,-1936260,-1936250,-1936239,-1936229,-1936218,-1936208,-1936197,-1936187,-1936176,-1936166,-1936155,-1936145,-1936134,-1936124,-1936113,-1936103,-1936092,-1936082,-1936071,-1936061,-1936050,-1936040,-1936029,-1936019,-1936008,-1935998,-1935987,-1935977,-1935966,-1935956,-1935945,-1935935,-1935924,-1935914,-1935903,-1935893,-1935882,-1935872,-1935861,-1935851,-1935840,-1935830,-1935819,-1935809,-1935798,-1935788,-1935777,-1935767,-1935756,-1935746,-1935735,-1935725,-1935714,-1935704,-1935693,-1935683,-1935672,-1935662,-1935651,-1935641,-1935630,-1935620,-1935609,-1935599,-1935588,-1935578,-1935567,-1935556,-1935546,-1935535,-1935525,-1935514,-1935504,-1935493,-1935483,-1935472,-1935462,-1935451,-1935441,-1935430,-1935420,-1935409,-1935399,-1935388,-1935378,-1935367,-1935357,-1935346,-1935336,-1935325,-1935315,-1935304,-1935293,-1935283,-1935272,-1935262,-1935251,-1935241,-1935230,-1935220,-1935209,-1935199,-1935188,-1935178,-1935167,-1935157,-1935146,-1935136,-1935125,-1935114,-1935104,-1935093,-1935083,-1935072,-1935062,-1935051,-1935041,-1935030,-1935020,-1935009,-1934999,-1934988,-1934978,-1934967,-1934956,-1934946,-1934935,-1934925,-1934914,-1934904,-1934893,-1934883,-1934872,-1934862,-1934851,-1934841,-1934830,-1934819,-1934809,-1934798,-1934788,-1934777,-1934767,-1934756,-1934746,-1934735,-1934725,-1934714,-1934703,-1934693,-1934682,-1934672,-1934661,-1934651,-1934640,-1934630,-1934619,-1934609,-1934598,-1934587,-1934577,-1934566,-1934556,-1934545,-1934535,-1934524,-1934514,-1934503,-1934492,-1934482,-1934471,-1934461,-1934450,-1934440,-1934429,-1934419,-1934408,-1934397,-1934387,-1934376,-1934366,-1934355,-1934345,-1934334,-1934324,-1934313,-1934302,-1934292,-1934281,-1934271,-1934260,-1934250,-1934239,-1934229,-1934218,-1934207,-1934197,-1934186,-1934176,-1934165,-1934155,-1934144,-1934133,-1934123,-1934112,-1934102,-1934091,-1934081,-1934070,-1934060,-1934049,-1934038,-1934028,-1934017,-1934007,-1933996,-1933986,-1933975,-1933964,-1933954,-1933943,-1933933,-1933922,-1933912,-1933901,-1933890,-1933880,-1933869,-1933859,-1933848,-1933838,-1933827,-1933816,-1933806,-1933795,-1933785,-1933774,-1933763,-1933753,-1933742,-1933732,-1933721,-1933711,-1933700,-1933689,-1933679,-1933668,-1933658,-1933647,-1933637,-1933626,-1933615,-1933605,-1933594,-1933584,-1933573,-1933562,-1933552,-1933541,-1933531,-1933520,-1933510,-1933499,-1933488,-1933478,-1933467,-1933457,-1933446,-1933435,-1933425,-1933414,-1933404,-1933393,-1933382,-1933372,-1933361,-1933351,-1933340,-1933330,-1933319,-1933308,-1933298,-1933287,-1933277,-1933266,-1933255,-1933245,-1933234,-1933224,-1933213,-1933202,-1933192,-1933181,-1933171,-1933160,-1933149,-1933139,-1933128,-1933118,-1933107,-1933096,-1933086,-1933075,-1933065,-1933054,-1933043,-1933033,-1933022,-1933012,-1933001,-1932990,-1932980,-1932969,-1932959,-1932948,-1932937,-1932927,-1932916,-1932906,-1932895,-1932884,-1932874,-1932863,-1932852,-1932842,-1932831,-1932821,-1932810,-1932799,-1932789,-1932778,-1932768,-1932757,-1932746,-1932736,-1932725,-1932715,-1932704,-1932693,-1932683,-1932672,-1932661,-1932651,-1932640,-1932630,-1932619,-1932608,-1932598,-1932587,-1932577,-1932566,-1932555,-1932545,-1932534,-1932523,-1932513,-1932502,-1932492,-1932481,-1932470,-1932460,-1932449,-1932438,-1932428,-1932417,-1932407,-1932396,-1932385,-1932375,-1932364,-1932353,-1932343,-1932332,-1932322,-1932311,-1932300,-1932290,-1932279,-1932268,-1932258,-1932247,-1932237,-1932226,-1932215,-1932205,-1932194,-1932183,-1932173,-1932162,-1932152,-1932141,-1932130,-1932120,-1932109,-1932098,-1932088,-1932077,-1932066,-1932056,-1932045,-1932035,-1932024,-1932013,-1932003,-1931992,-1931981,-1931971,-1931960,-1931949,-1931939,-1931928,-1931918,-1931907,-1931896,-1931886,-1931875,-1931864,-1931854,-1931843,-1931832,-1931822,-1931811,-1931800,-1931790,-1931779,-1931769,-1931758,-1931747,-1931737,-1931726,-1931715,-1931705,-1931694,-1931683,-1931673,-1931662,-1931651,-1931641,-1931630,-1931619,-1931609,-1931598,-1931588,-1931577,-1931566,-1931556,-1931545,-1931534,-1931524,-1931513,-1931502,-1931492,-1931481,-1931470,-1931460,-1931449,-1931438,-1931428,-1931417,-1931406,-1931396,-1931385,-1931374,-1931364,-1931353,-1931342,-1931332,-1931321,-1931310,-1931300,-1931289,-1931278,-1931268,-1931257,-1931247,-1931236,-1931225,-1931215,-1931204,-1931193,-1931183,-1931172,-1931161,-1931151,-1931140,-1931129,-1931119,-1931108,-1931097,-1931087,-1931076,-1931065,-1931055,-1931044,-1931033,-1931023,-1931012,-1931001,-1930990,-1930980,-1930969,-1930958,-1930948,-1930937,-1930926,-1930916,-1930905,-1930894,-1930884,-1930873,-1930862,-1930852,-1930841,-1930830,-1930820,-1930809,-1930798,-1930788,-1930777,-1930766,-1930756,-1930745,-1930734,-1930724,-1930713,-1930702,-1930692,-1930681,-1930670,-1930660,-1930649,-1930638,-1930627,-1930617,-1930606,-1930595,-1930585,-1930574,-1930563,-1930553,-1930542,-1930531,-1930521,-1930510,-1930499,-1930489,-1930478,-1930467,-1930456,-1930446,-1930435,-1930424,-1930414,-1930403,-1930392,-1930382,-1930371,-1930360,-1930350,-1930339,-1930328,-1930317,-1930307,-1930296,-1930285,-1930275,-1930264,-1930253,-1930243,-1930232,-1930221,-1930211,-1930200,-1930189,-1930178,-1930168,-1930157,-1930146,-1930136,-1930125,-1930114,-1930104,-1930093,-1930082,-1930071,-1930061,-1930050,-1930039,-1930029,-1930018,-1930007,-1929997,-1929986,-1929975,-1929964,-1929954,-1929943,-1929932,-1929922,-1929911,-1929900,-1929889,-1929879,-1929868,-1929857,-1929847,-1929836,-1929825,-1929814,-1929804,-1929793,-1929782,-1929772,-1929761,-1929750,-1929739,-1929729,-1929718,-1929707,-1929697,-1929686,-1929675,-1929664,-1929654,-1929643,-1929632,-1929622,-1929611,-1929600,-1929589,-1929579,-1929568,-1929557,-1929547,-1929536,-1929525,-1929514,-1929504,-1929493,-1929482,-1929472,-1929461,-1929450,-1929439,-1929429,-1929418,-1929407,-1929396,-1929386,-1929375,-1929364,-1929354,-1929343,-1929332,-1929321,-1929311,-1929300,-1929289,-1929278,-1929268,-1929257,-1929246,-1929236,-1929225,-1929214,-1929203,-1929193,-1929182,-1929171,-1929160,-1929150,-1929139,-1929128,-1929118,-1929107,-1929096,-1929085,-1929075,-1929064,-1929053,-1929042,-1929032,-1929021,-1929010,-1928999,-1928989,-1928978,-1928967,-1928956,-1928946,-1928935,-1928924,-1928914,-1928903,-1928892,-1928881,-1928871,-1928860,-1928849,-1928838,-1928828,-1928817,-1928806,-1928795,-1928785,-1928774,-1928763,-1928752,-1928742,-1928731,-1928720,-1928709,-1928699,-1928688,-1928677,-1928666,-1928656,-1928645,-1928634,-1928623,-1928613,-1928602,-1928591,-1928580,-1928570,-1928559,-1928548,-1928537,-1928527,-1928516,-1928505,-1928494,-1928484,-1928473,-1928462,-1928451,-1928441,-1928430,-1928419,-1928408,-1928398,-1928387,-1928376,-1928365,-1928354,-1928344,-1928333,-1928322,-1928311,-1928301,-1928290,-1928279,-1928268,-1928258,-1928247,-1928236,-1928225,-1928215,-1928204,-1928193,-1928182,-1928172,-1928161,-1928150,-1928139,-1928128,-1928118,-1928107,-1928096,-1928085,-1928075,-1928064,-1928053,-1928042,-1928032,-1928021,-1928010,-1927999,-1927988,-1927978,-1927967,-1927956,-1927945,-1927935,-1927924,-1927913,-1927902,-1927891,-1927881,-1927870,-1927859,-1927848,-1927838,-1927827,-1927816,-1927805,-1927795,-1927784,-1927773,-1927762,-1927751,-1927741,-1927730,-1927719,-1927708,-1927697,-1927687,-1927676,-1927665,-1927654,-1927644,-1927633,-1927622,-1927611,-1927600,-1927590,-1927579,-1927568,-1927557,-1927547,-1927536,-1927525,-1927514,-1927503,-1927493,-1927482,-1927471,-1927460,-1927449,-1927439,-1927428,-1927417,-1927406,-1927395,-1927385,-1927374,-1927363,-1927352,-1927342,-1927331,-1927320,-1927309,-1927298,-1927288,-1927277,-1927266,-1927255,-1927244,-1927234,-1927223,-1927212,-1927201,-1927190,-1927180,-1927169,-1927158,-1927147,-1927136,-1927126,-1927115,-1927104,-1927093,-1927082,-1927072,-1927061,-1927050,-1927039,-1927028,-1927018,-1927007,-1926996,-1926985,-1926974,-1926964,-1926953,-1926942,-1926931,-1926920,-1926909,-1926899,-1926888,-1926877,-1926866,-1926855,-1926845,-1926834,-1926823,-1926812,-1926801,-1926791,-1926780,-1926769,-1926758,-1926747,-1926737,-1926726,-1926715,-1926704,-1926693,-1926682,-1926672,-1926661,-1926650,-1926639,-1926628,-1926618,-1926607,-1926596,-1926585,-1926574,-1926563,-1926553,-1926542,-1926531,-1926520,-1926509,-1926499,-1926488,-1926477,-1926466,-1926455,-1926444,-1926434,-1926423,-1926412,-1926401,-1926390,-1926379,-1926369,-1926358,-1926347,-1926336,-1926325,-1926315,-1926304,-1926293,-1926282,-1926271,-1926260,-1926250,-1926239,-1926228,-1926217,-1926206,-1926195,-1926185,-1926174,-1926163,-1926152,-1926141,-1926130,-1926120,-1926109,-1926098,-1926087,-1926076,-1926065,-1926055,-1926044,-1926033,-1926022,-1926011,-1926000,-1925990,-1925979,-1925968,-1925957,-1925946,-1925935,-1925925,-1925914,-1925903,-1925892,-1925881,-1925870,-1925859,-1925849,-1925838,-1925827,-1925816,-1925805,-1925794,-1925784,-1925773,-1925762,-1925751,-1925740,-1925729,-1925718,-1925708,-1925697,-1925686,-1925675,-1925664,-1925653,-1925643,-1925632,-1925621,-1925610,-1925599,-1925588,-1925577,-1925567,-1925556,-1925545,-1925534,-1925523,-1925512,-1925501,-1925491,-1925480,-1925469,-1925458,-1925447,-1925436,-1925425,-1925415,-1925404,-1925393,-1925382,-1925371,-1925360,-1925349,-1925339,-1925328,-1925317,-1925306,-1925295,-1925284,-1925273,-1925263,-1925252,-1925241,-1925230,-1925219,-1925208,-1925197,-1925187,-1925176,-1925165,-1925154,-1925143,-1925132,-1925121,-1925110,-1925100,-1925089,-1925078,-1925067,-1925056,-1925045,-1925034,-1925024,-1925013,-1925002,-1924991,-1924980,-1924969,-1924958,-1924947
);
signal constA1 : signed(w_coef-1 downto 0):= to_signed(A1(0),w_coef);

signal BP_out : signed(W_in-1 downto 0) := (others =>'0');
signal data_out_temp:  signed(W_in-1 downto 0) := (others =>'0');
signal BW_clk : std_logic := '0';
begin

process(CLK_50,nReset) 
variable counter : integer := 0;
variable direction: std_logic := '0';
begin
if (nReset = '0') then
	counter := 0;
	direction:= '0';
elsif (rising_edge(CLK_50)) then
	if (new_val = '1') then
	if (direction = '0') then
		constA1 <= to_signed(A1(counter),w_coef);
		counter := counter + 1;
		if(counter = Arr_size) then
			direction := '1';
		end if;
	end if;
	if(direction = '1') then
		counter := counter -1;
		constA1 <= to_signed(A1(counter),w_coef);
		if(counter = 0) then
			direction := '0';
		end if;
	end if;
	end if;
end if;
end process;

IIRDF_inst : IIRDF1_BW 
generic map(
   W_in => W_in,
	W_coef => W_coef,
	A0 => A0,
	A2 => A2,
	B0 => B0,
	B1 => B1,
	B2 => B2
)
port map(
	iCLK => CLK_50,          
	iRESET_N => nReset,      
	new_val => new_val,        
	IIR_in => data_in,                 
	IIR_out => BP_out,         
   A1 => constA1
);

process(CLK_50,nReset)
begin
if nReset = '0' then
	data_out <= (others => '0');
elsif(rising_edge(CLK_50)) then
	if(new_val = '1') then
	if WahWah_EN = '0' then
		data_out <= data_in;
	elsif WahWah_EN = '1' then
		data_out <= BP_out + data_in;
	end if;
	end if;
end if;
end process;
end;