library IEEE;
use IEEE.STD_LOGIC_1164.ALL;  
use IEEE.NUMERIC_STD.ALL;
use work.data_types.all;

entity impulsebench is
end;

architecture testbench of impulsebench is

	signal rst : std_logic := '0';
	signal clk : std_logic := '0';
	signal interclk : std_logic := '0';
	signal sndclk : std_logic := '0';
	signal word : signed(15 downto 0);
	signal inter : signed(15 downto 0);
  signal resp : signed(15 downto 0);

  component polyphase
    Generic (
        coef_scale : integer;
        w_acc : integer;
        coef : array_of_integers;
        D : integer
    );
    port (
      rst    : in std_logic;
      clk    : in std_logic;
      inclk : in std_logic;
      outclk : out std_logic;
      word   : in signed(15 downto 0);
      resp   : out signed(15 downto 0)
    );
  end component;

    
begin
  rst <= '1' AFTER 20 ns; -- reset pin
  clk <= NOT clk AFTER 10 ns; -- "fast clock"; 50 MHz klok

  process(clk)
    variable counter: integer := 0;
  begin
    if rising_edge(clk) then
      counter := counter + 1;
      if counter < 3000 then
        word <= x"0000";
      elsif counter < 100000 then
        word <= x"3fff";
      else
        word <= -word;
      end if;
    end if;
  end process;

  filter_inst1 : polyphase
  generic map (
    coef_scale => 2**16,
    w_acc => 32,
    D => 64,
    coef => (
-10,-9,-20,-36,-52,-65,-64,-40,15,108,239,399,575,745,886,978,1008,970,870,724,553,378,221,94,6,-45,-65,-64,-50,-34,-19,-8,
-4,-10,-22,-38,-54,-65,-62,-35,25,123,258,421,597,764,900,986,1007,961,854,704,531,357,203,81,-2,-49,-66,-62,-48,-32,-17,-7,
-4,-12,-24,-40,-56,-66,-60,-30,35,138,277,443,619,783,914,992,1005,950,838,683,509,337,186,69,-10,-52,-66,-61,-46,-30,-16,-6,
-5,-13,-26,-42,-58,-66,-58,-24,45,153,296,464,640,802,927,997,1001,939,820,662,486,316,169,57,-17,-56,-66,-59,-44,-28,-14,-6,
-6,-14,-28,-44,-59,-66,-56,-17,57,169,316,486,662,820,939,1001,997,927,802,640,464,296,153,45,-24,-58,-66,-58,-42,-26,-13,-5,
-6,-16,-30,-46,-61,-66,-52,-10,69,186,337,509,683,838,950,1005,992,914,783,619,443,277,138,35,-30,-60,-66,-56,-40,-24,-12,-4,
-7,-17,-32,-48,-62,-66,-49,-2,81,203,357,531,704,854,961,1007,986,900,764,597,421,258,123,25,-35,-62,-65,-54,-38,-22,-10,-4,
-8,-19,-34,-50,-64,-65,-45,6,94,221,378,553,724,870,970,1008,978,886,745,575,399,239,108,15,-40,-64,-65,-52,-36,-20,-9,-10
  )
  )
  port map (
    rst => rst,
    clk => clk,
    inclk => clk,
    outclk => interclk,
    word => word,
    resp => inter
  );
  filter_inst2 : polyphase
  generic map (
    coef_scale => 2**16,
    w_acc => 32,
    D => 16,
    coef => (
-0,0,-0,-1,-3,-4,-2,6,21,36,40,13,-56,-167,-300,-435,3672,-332,-280,-176,-73,-1,32,35,22,8,-1,-3,-2,-1,-0,0,
0,0,-0,-1,-3,-4,-4,3,18,37,47,28,-37,-153,-311,-530,3634,-226,-252,-180,-88,-15,24,32,23,10,1,-2,-2,-1,-0,-0,
0,0,0,-1,-3,-5,-5,1,16,37,52,42,-16,-133,-313,-615,3558,-119,-217,-177,-99,-28,15,28,23,11,2,-2,-2,-1,-0,-0,
0,0,0,-1,-2,-5,-6,-2,12,35,56,54,6,-108,-305,-687,3447,-15,-177,-170,-107,-40,5,24,22,12,4,-1,-2,-1,-0,-0,
0,0,0,-0,-2,-5,-8,-5,8,32,58,66,29,-80,-287,-742,3302,83,-133,-157,-112,-51,-4,19,21,13,5,-0,-1,-1,-0,-0,
0,0,0,-0,-2,-5,-9,-7,4,28,59,76,51,-48,-260,-777,3126,174,-86,-140,-113,-60,-13,13,19,13,6,1,-1,-1,-0,-0,
0,0,0,0,-2,-5,-9,-10,-0,24,57,83,72,-13,-223,-789,2921,254,-38,-119,-111,-66,-21,7,16,13,6,1,-1,-1,-0,-0,
0,0,0,0,-1,-5,-10,-12,-5,18,54,88,91,23,-177,-778,2693,322,9,-95,-105,-71,-28,1,13,13,7,2,-0,-1,-0,-0,
0,0,1,1,-1,-4,-10,-14,-9,11,49,91,108,59,-124,-740,2445,377,55,-69,-96,-73,-35,-4,10,12,7,3,0,-1,-0,-0,
0,0,1,1,-0,-4,-10,-16,-14,4,42,90,122,94,-65,-674,2181,418,97,-41,-84,-73,-40,-10,7,10,7,3,0,-0,-0,-0,
0,0,1,1,0,-3,-9,-17,-18,-3,34,87,133,128,-2,-581,1906,444,135,-13,-70,-70,-44,-15,3,9,7,3,1,-0,-0,-0,
0,0,1,1,1,-2,-9,-17,-22,-10,24,81,139,158,65,-459,1625,455,168,15,-55,-66,-46,-19,-0,7,7,4,1,-0,-0,-0,
0,0,1,1,2,-1,-8,-18,-25,-18,14,72,142,185,132,-309,1343,452,195,42,-38,-60,-47,-23,-4,5,6,4,1,0,-0,-0,
-0,0,1,2,2,0,-6,-17,-27,-25,3,61,140,206,198,-133,1064,436,215,67,-20,-51,-46,-26,-7,3,5,4,1,0,-0,-0,
-0,0,1,2,3,1,-5,-16,-29,-31,-9,48,133,221,260,68,793,407,227,89,-2,-42,-44,-28,-10,1,5,4,2,0,-0,-0,
-0,0,1,2,3,2,-3,-15,-29,-36,-20,32,122,230,317,291,534,367,232,107,16,-32,-41,-29,-12,-1,4,3,2,0,0,-0,
-0,0,0,2,3,4,-1,-12,-29,-41,-32,16,107,232,367,534,291,317,230,122,32,-20,-36,-29,-15,-3,2,3,2,1,0,-0,
-0,-0,0,2,4,5,1,-10,-28,-44,-42,-2,89,227,407,793,68,260,221,133,48,-9,-31,-29,-16,-5,1,3,2,1,0,-0,
-0,-0,0,1,4,5,3,-7,-26,-46,-51,-20,67,215,436,1064,-133,198,206,140,61,3,-25,-27,-17,-6,0,2,2,1,0,-0,
-0,-0,0,1,4,6,5,-4,-23,-47,-60,-38,42,195,452,1343,-309,132,185,142,72,14,-18,-25,-18,-8,-1,2,1,1,0,0,
-0,-0,-0,1,4,7,7,-0,-19,-46,-66,-55,15,168,455,1625,-459,65,158,139,81,24,-10,-22,-17,-9,-2,1,1,1,0,0,
-0,-0,-0,1,3,7,9,3,-15,-44,-70,-70,-13,135,444,1906,-581,-2,128,133,87,34,-3,-18,-17,-9,-3,0,1,1,0,0,
-0,-0,-0,0,3,7,10,7,-10,-40,-73,-84,-41,97,418,2181,-674,-65,94,122,90,42,4,-14,-16,-10,-4,-0,1,1,0,0,
-0,-0,-1,0,3,7,12,10,-4,-35,-73,-96,-69,55,377,2445,-740,-124,59,108,91,49,11,-9,-14,-10,-4,-1,1,1,0,0,
-0,-0,-1,-0,2,7,13,13,1,-28,-71,-105,-95,9,322,2693,-778,-177,23,91,88,54,18,-5,-12,-10,-5,-1,0,0,0,0,
-0,-0,-1,-1,1,6,13,16,7,-21,-66,-111,-119,-38,254,2921,-789,-223,-13,72,83,57,24,-0,-10,-9,-5,-2,0,0,0,0,
-0,-0,-1,-1,1,6,13,19,13,-13,-60,-113,-140,-86,174,3126,-777,-260,-48,51,76,59,28,4,-7,-9,-5,-2,-0,0,0,0,
-0,-0,-1,-1,-0,5,13,21,19,-4,-51,-112,-157,-133,83,3302,-742,-287,-80,29,66,58,32,8,-5,-8,-5,-2,-0,0,0,0,
-0,-0,-1,-2,-1,4,12,22,24,5,-40,-107,-170,-177,-15,3447,-687,-305,-108,6,54,56,35,12,-2,-6,-5,-2,-1,0,0,0,
-0,-0,-1,-2,-2,2,11,23,28,15,-28,-99,-177,-217,-119,3558,-615,-313,-133,-16,42,52,37,16,1,-5,-5,-3,-1,0,0,0,
-0,-0,-1,-2,-2,1,10,23,32,24,-15,-88,-180,-252,-226,3634,-530,-311,-153,-37,28,47,37,18,3,-4,-4,-3,-1,-0,0,0,
0,-0,-1,-2,-3,-1,8,22,35,32,-1,-73,-176,-280,-332,3672,-435,-300,-167,-56,13,40,36,21,6,-2,-4,-3,-1,-0,0,-0
  )
  )
  port map (
    rst => rst,
    clk => clk,
    inclk => interclk,
    outclk => sndclk,
    word => inter,
    resp => resp
  );
end;
