library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity WahWah_FX is
port (
	CLK_50		: in std_logic;
	nReset		: in std_logic;
	new_val		: in std_logic;       -- indicates a new input value, input from data_over
	data_in		: in signed (15 downto 0);         
	data_out		: out signed (15 downto 0);   -- Output
	WahWah_EN 	: in std_logic
);
end entity WahWah_FX;

architecture behaviour of WahWah_FX is
constant W_coef : integer := 23;
constant W_in : integer := 16;
constant A0 : integer :=1048576 ;
constant A2 : integer :=1034939 ;
constant B0 : integer :=6818 ;
constant B1 : integer := 0;
constant B2 : integer := -6818 ; 
constant Arr_size : integer := 1250;

component IIRDF1_BW is
generic (
   W_in : integer ;
	W_coef : integer;
	A0 : integer;
	A2 : integer;
	B0 : integer ;
	B1 : integer;
	B2 : integer    
);
port (
	iCLK            : in std_logic;
	iRESET_N        : in std_logic;
	new_val         : in std_logic;       -- indicates a new input value, input from data_over
	IIR_in          : in signed (15 downto 0);   -- singed is expected             
	IIR_out         : out signed (15 downto 0);   -- Output
   A1 : in signed(W_coef-1 downto 0)

);
end component;


type cA1_array_type is array (0 to Arr_size) of integer;
signal A1 : cA1_array_type:=(-2079063,-2079027,-2078991,-2078955,-2078919,-2078882,-2078846,-2078809,-2078772,-2078735,-2078698,-2078660,-2078623,-2078585,-2078548,-2078510,-2078472,-2078434,-2078395,-2078357,-2078318,-2078279,-2078241,-2078202,-2078162,-2078123,-2078084,-2078044,-2078004,-2077964,-2077924,-2077884,-2077844,-2077803,-2077763,-2077722,-2077681,-2077640,-2077599,-2077558,-2077516,-2077475,-2077433,-2077391,-2077349,-2077307,-2077265,-2077222,-2077180,-2077137,-2077094,-2077051,-2077008,-2076965,-2076921,-2076878,-2076834,-2076790,-2076746,-2076702,-2076658,-2076613,-2076569,-2076524,-2076479,-2076434,-2076389,-2076344,-2076298,-2076253,-2076207,-2076161,-2076115,-2076069,-2076023,-2075976,-2075930,-2075883,-2075836,-2075789,-2075742,-2075695,-2075647,-2075600,-2075552,-2075504,-2075456,-2075408,-2075360,-2075311,-2075263,-2075214,-2075165,-2075116,-2075067,-2075018,-2074968,-2074919,-2074869,-2074819,-2074769,-2074719,-2074669,-2074618,-2074568,-2074517,-2074466,-2074415,-2074364,-2074313,-2074262,-2074210,-2074158,-2074106,-2074054,-2074002,-2073950,-2073898,-2073845,-2073792,-2073740,-2073687,-2073634,-2073580,-2073527,-2073473,-2073420,-2073366,-2073312,-2073258,-2073204,-2073149,-2073095,-2073040,-2072985,-2072930,-2072875,-2072820,-2072764,-2072709,-2072653,-2072597,-2072542,-2072485,-2072429,-2072373,-2072316,-2072260,-2072203,-2072146,-2072089,-2072032,-2071974,-2071917,-2071859,-2071801,-2071743,-2071685,-2071627,-2071569,-2071510,-2071451,-2071393,-2071334,-2071275,-2071215,-2071156,-2071097,-2071037,-2070977,-2070917,-2070857,-2070797,-2070737,-2070676,-2070615,-2070555,-2070494,-2070433,-2070371,-2070310,-2070249,-2070187,-2070125,-2070063,-2070001,-2069939,-2069877,-2069814,-2069752,-2069689,-2069626,-2069563,-2069500,-2069436,-2069373,-2069309,-2069246,-2069182,-2069118,-2069053,-2068989,-2068925,-2068860,-2068795,-2068730,-2068665,-2068600,-2068535,-2068469,-2068404,-2068338,-2068272,-2068206,-2068140,-2068074,-2068007,-2067941,-2067874,-2067807,-2067740,-2067673,-2067605,-2067538,-2067470,-2067403,-2067335,-2067267,-2067199,-2067130,-2067062,-2066993,-2066925,-2066856,-2066787,-2066718,-2066648,-2066579,-2066509,-2066440,-2066370,-2066300,-2066230,-2066159,-2066089,-2066018,-2065948,-2065877,-2065806,-2065735,-2065663,-2065592,-2065520,-2065449,-2065377,-2065305,-2065233,-2065161,-2065088,-2065016,-2064943,-2064870,-2064797,-2064724,-2064651,-2064577,-2064504,-2064430,-2064356,-2064282,-2064208,-2064134,-2064060,-2063985,-2063911,-2063836,-2063761,-2063686,-2063610,-2063535,-2063460,-2063384,-2063308,-2063232,-2063156,-2063080,-2063003,-2062927,-2062850,-2062774,-2062697,-2062620,-2062542,-2062465,-2062387,-2062310,-2062232,-2062154,-2062076,-2061998,-2061920,-2061841,-2061762,-2061684,-2061605,-2061526,-2061447,-2061367,-2061288,-2061208,-2061128,-2061048,-2060968,-2060888,-2060808,-2060727,-2060647,-2060566,-2060485,-2060404,-2060323,-2060242,-2060160,-2060079,-2059997,-2059915,-2059833,-2059751,-2059669,-2059586,-2059504,-2059421,-2059338,-2059255,-2059172,-2059089,-2059005,-2058922,-2058838,-2058754,-2058670,-2058586,-2058502,-2058417,-2058333,-2058248,-2058163,-2058078,-2057993,-2057908,-2057822,-2057737,-2057651,-2057565,-2057479,-2057393,-2057307,-2057221,-2057134,-2057047,-2056961,-2056874,-2056787,-2056699,-2056612,-2056524,-2056437,-2056349,-2056261,-2056173,-2056085,-2055996,-2055908,-2055819,-2055730,-2055642,-2055552,-2055463,-2055374,-2055284,-2055195,-2055105,-2055015,-2054925,-2054835,-2054745,-2054654,-2054563,-2054473,-2054382,-2054291,-2054200,-2054108,-2054017,-2053925,-2053833,-2053742,-2053650,-2053557,-2053465,-2053373,-2053280,-2053187,-2053094,-2053001,-2052908,-2052815,-2052722,-2052628,-2052534,-2052440,-2052346,-2052252,-2052158,-2052064,-2051969,-2051874,-2051779,-2051685,-2051589,-2051494,-2051399,-2051303,-2051208,-2051112,-2051016,-2050920,-2050823,-2050727,-2050630,-2050534,-2050437,-2050340,-2050243,-2050146,-2050048,-2049951,-2049853,-2049755,-2049657,-2049559,-2049461,-2049363,-2049264,-2049166,-2049067,-2048968,-2048869,-2048770,-2048670,-2048571,-2048471,-2048372,-2048272,-2048172,-2048071,-2047971,-2047871,-2047770,-2047669,-2047569,-2047467,-2047366,-2047265,-2047164,-2047062,-2046960,-2046858,-2046756,-2046654,-2046552,-2046450,-2046347,-2046244,-2046141,-2046038,-2045935,-2045832,-2045729,-2045625,-2045521,-2045418,-2045314,-2045210,-2045105,-2045001,-2044896,-2044792,-2044687,-2044582,-2044477,-2044372,-2044266,-2044161,-2044055,-2043949,-2043843,-2043737,-2043631,-2043525,-2043418,-2043312,-2043205,-2043098,-2042991,-2042884,-2042776,-2042669,-2042561,-2042454,-2042346,-2042238,-2042130,-2042021,-2041913,-2041804,-2041696,-2041587,-2041478,-2041368,-2041259,-2041150,-2041040,-2040931,-2040821,-2040711,-2040601,-2040490,-2040380,-2040269,-2040159,-2040048,-2039937,-2039826,-2039715,-2039603,-2039492,-2039380,-2039268,-2039156,-2039044,-2038932,-2038820,-2038707,-2038594,-2038482,-2038369,-2038256,-2038142,-2038029,-2037916,-2037802,-2037688,-2037574,-2037460,-2037346,-2037232,-2037117,-2037003,-2036888,-2036773,-2036658,-2036543,-2036428,-2036312,-2036197,-2036081,-2035965,-2035849,-2035733,-2035617,-2035500,-2035384,-2035267,-2035150,-2035033,-2034916,-2034799,-2034681,-2034564,-2034446,-2034328,-2034211,-2034092,-2033974,-2033856,-2033737,-2033619,-2033500,-2033381,-2033262,-2033143,-2033023,-2032904,-2032784,-2032665,-2032545,-2032425,-2032304,-2032184,-2032064,-2031943,-2031822,-2031701,-2031580,-2031459,-2031338,-2031217,-2031095,-2030973,-2030851,-2030729,-2030607,-2030485,-2030363,-2030240,-2030117,-2029995,-2029872,-2029749,-2029625,-2029502,-2029378,-2029255,-2029131,-2029007,-2028883,-2028759,-2028634,-2028510,-2028385,-2028261,-2028136,-2028011,-2027885,-2027760,-2027635,-2027509,-2027383,-2027257,-2027131,-2027005,-2026879,-2026752,-2026626,-2026499,-2026372,-2026245,-2026118,-2025991,-2025864,-2025736,-2025608,-2025480,-2025353,-2025224,-2025096,-2024968,-2024839,-2024711,-2024582,-2024453,-2024324,-2024195,-2024065,-2023936,-2023806,-2023676,-2023546,-2023416,-2023286,-2023156,-2023025,-2022895,-2022764,-2022633,-2022502,-2022371,-2022240,-2022108,-2021977,-2021845,-2021713,-2021581,-2021449,-2021317,-2021184,-2021052,-2020919,-2020786,-2020653,-2020520,-2020387,-2020254,-2020120,-2019987,-2019853,-2019719,-2019585,-2019451,-2019316,-2019182,-2019047,-2018912,-2018778,-2018643,-2018507,-2018372,-2018237,-2018101,-2017965,-2017829,-2017693,-2017557,-2017421,-2017285,-2017148,-2017011,-2016875,-2016738,-2016600,-2016463,-2016326,-2016188,-2016051,-2015913,-2015775,-2015637,-2015499,-2015360,-2015222,-2015083,-2014944,-2014805,-2014666,-2014527,-2014388,-2014248,-2014109,-2013969,-2013829,-2013689,-2013549,-2013409,-2013268,-2013128,-2012987,-2012846,-2012705,-2012564,-2012423,-2012282,-2012140,-2011998,-2011857,-2011715,-2011573,-2011430,-2011288,-2011146,-2011003,-2010860,-2010717,-2010574,-2010431,-2010288,-2010144,-2010001,-2009857,-2009713,-2009569,-2009425,-2009281,-2009136,-2008992,-2008847,-2008702,-2008557,-2008412,-2008267,-2008121,-2007976,-2007830,-2007685,-2007539,-2007393,-2007246,-2007100,-2006953,-2006807,-2006660,-2006513,-2006366,-2006219,-2006072,-2005924,-2005777,-2005629,-2005481,-2005333,-2005185,-2005037,-2004888,-2004740,-2004591,-2004442,-2004293,-2004144,-2003995,-2003846,-2003696,-2003546,-2003397,-2003247,-2003097,-2002946,-2002796,-2002646,-2002495,-2002344,-2002193,-2002042,-2001891,-2001740,-2001589,-2001437,-2001285,-2001133,-2000981,-2000829,-2000677,-2000525,-2000372,-2000220,-2000067,-1999914,-1999761,-1999608,-1999454,-1999301,-1999147,-1998993,-1998839,-1998685,-1998531,-1998377,-1998222,-1998068,-1997913,-1997758,-1997603,-1997448,-1997293,-1997138,-1996982,-1996826,-1996670,-1996515,-1996358,-1996202,-1996046,-1995889,-1995733,-1995576,-1995419,-1995262,-1995105,-1994948,-1994790,-1994632,-1994475,-1994317,-1994159,-1994001,-1993842,-1993684,-1993526,-1993367,-1993208,-1993049,-1992890,-1992731,-1992571,-1992412,-1992252,-1992092,-1991933,-1991772,-1991612,-1991452,-1991291,-1991131,-1990970,-1990809,-1990648,-1990487,-1990326,-1990164,-1990003,-1989841,-1989679,-1989517,-1989355,-1989193,-1989031,-1988868,-1988706,-1988543,-1988380,-1988217,-1988054,-1987890,-1987727,-1987563,-1987400,-1987236,-1987072,-1986908,-1986743,-1986579,-1986414,-1986250,-1986085,-1985920,-1985755,-1985589,-1985424,-1985259,-1985093,-1984927,-1984761,-1984595,-1984429,-1984263,-1984096,-1983930,-1983763,-1983596,-1983429,-1983262,-1983095,-1982927,-1982760,-1982592,-1982424,-1982256,-1982088,-1981920,-1981752,-1981583,-1981415,-1981246,-1981077,-1980908,-1980739,-1980569,-1980400,-1980230,-1980061,-1979891,-1979721,-1979551,-1979380,-1979210,-1979039,-1978869,-1978698,-1978527,-1978356,-1978185,-1978013,-1977842,-1977670,-1977499,-1977327,-1977155,-1976983,-1976810,-1976638,-1976465,-1976293,-1976120,-1975947,-1975774,-1975600,-1975427,-1975254,-1975080,-1974906,-1974732,-1974558,-1974384,-1974210,-1974035,-1973861,-1973686,-1973511,-1973336,-1973161,-1972986,-1972810,-1972635,-1972459,-1972283,-1972107,-1971931,-1971755,-1971579,-1971402,-1971225,-1971049,-1970872,-1970695,-1970518,-1970340,-1970163,-1969985,-1969808,-1969630,-1969452,-1969274,-1969095,-1968917,-1968739,-1968560,-1968381,-1968202,-1968023,-1967844,-1967665,-1967485,-1967306,-1967126,-1966946,-1966766,-1966586,-1966406,-1966225,-1966045,-1965864,-1965683,-1965502,-1965321,-1965140,-1964959,-1964777,-1964596,-1964414,-1964232,-1964050,-1963868,-1963686,-1963503,-1963321,-1963138,-1962955,-1962772,-1962589,-1962406,-1962222,-1962039,-1961855,-1961672,-1961488,-1961304,-1961119,-1960935,-1960751,-1960566,-1960381,-1960197,-1960012,-1959826,-1959641,-1959456,-1959270,-1959085,-1958899,-1958713,-1958527,-1958341,-1958154,-1957968,-1957781,-1957595,-1957408,-1957221,-1957034,-1956846,-1956659,-1956472,-1956284,-1956096,-1955908,-1955720,-1955532,-1955344,-1955155,-1954967,-1954778,-1954589,-1954400,-1954211,-1954022,-1953832,-1953643,-1953453,-1953263,-1953073,-1952883,-1952693,-1952503,-1952312,-1952122,-1951931,-1951740,-1951549,-1951358,-1951166,-1950975,-1950784,-1950592,-1950400,-1950208,-1950016,-1949824,-1949631,-1949439,-1949246,-1949054,-1948861,-1948668,-1948475,-1948281,-1948088,-1947894,-1947701,-1947507,-1947313,-1947119,-1946925,-1946730,-1946536,-1946341,-1946146,-1945952,-1945757,-1945561,-1945366,-1945171,-1944975,-1944779,-1944584,-1944388,-1944192,-1943995,-1943799,-1943603,-1943406,-1943209,-1943012,-1942815,-1942618,-1942421,-1942223,-1942026,-1941828,-1941630,-1941433,-1941234,-1941036,-1940838,-1940639,-1940441,-1940242,-1940043,-1939844,-1939645,-1939446,-1939246,-1939047,-1938847,-1938647,-1938447,-1938247,-1938047,-1937847,-1937646,-1937446,-1937245,-1937044,-1936843,-1936642,-1936441,-1936239,-1936038,-1935836,-1935634,-1935432,-1935230,-1935028,-1934826,-1934623,-1934421,-1934218,-1934015,-1933812,-1933609,-1933406,-1933202,-1932999,-1932795,-1932591,-1932387,-1932183,-1931979,-1931775,-1931570,-1931366,-1931161,-1930956,-1930751,-1930546,-1930341,-1930136,-1929930,-1929724,-1929519,-1929313,-1929107,-1928901,-1928694,-1928488,-1928281,-1928075,-1927868,-1927661,-1927454,-1927247,-1927039,-1926832,-1926624,-1926416,-1926208,-1926000,-1925792,-1925584,-1925376,-1925167,-1924958,-1924749
);
signal constA1 : signed(w_coef-1 downto 0):= to_signed(A1(0),w_coef);

signal BP_out : signed(W_in-1 downto 0) := (others =>'0');
signal data_out_temp:  signed(W_in-1 downto 0) := (others =>'0');
signal BW_clk : std_logic := '0';
begin

process(CLK_50,nReset) 
variable counter : integer := 0;
variable direction: std_logic := '0';
begin
if (nReset = '0') then
	counter := 0;
	direction:= '0';
elsif (rising_edge(CLK_50)) then
	if (new_val = '1') then
	if (direction = '0') then
		constA1 <= to_signed(A1(counter),w_coef);
		counter := counter + 1;
		if(counter = Arr_size) then
			direction := '1';
		end if;
	end if;
	if(direction = '1') then
		counter := counter -1;
		constA1 <= to_signed(A1(counter),w_coef);
		if(counter = 0) then
			direction := '0';
		end if;
	end if;
	end if;
end if;
end process;

IIRDF_inst : IIRDF1_BW 
generic map(
   W_in => W_in,
	W_coef => W_coef,
	A0 => A0,
	A2 => A2,
	B0 => B0,
	B1 => B1,
	B2 => B2
)
port map(
	iCLK => CLK_50,          
	iRESET_N => nReset,      
	new_val => new_val,        
	IIR_in => data_in,                 
	IIR_out => BP_out,         
   A1 => constA1
);

process(CLK_50,nReset)
begin
if nReset = '0' then
	data_out <= (others => '0');
elsif(rising_edge(CLK_50)) then
	if(new_val = '1') then
	if WahWah_EN = '0' then
		data_out <= data_in;
	elsif WahWah_EN = '1' then
		data_out <= BP_out + data_in;
	end if;
	end if;
end if;
end process;
end;