library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity WahWah_FX is
port (
	CLK_50		: in std_logic;
	nReset		: in std_logic;
	new_val		: in std_logic;       -- indicates a new input value, input from data_over
	data_in		: in signed (15 downto 0);         
	data_out		: out signed (15 downto 0);   -- Output
	WahWah_EN 	: in std_logic
);
end entity WahWah_FX;

architecture behaviour of WahWah_FX is
constant W_coef : integer := 20;
constant W_in : integer := 16;


component IIRDF1 is
generic (
    W_in : integer ;
	 W_coef : integer   
);
port (
	iCLK            : in std_logic;
	iRESET_N        : in std_logic;
	new_val         : in std_logic;       -- indicates a new input value, input from data_over
	IIR_in          : in signed (15 downto 0);   -- singed is expected             
	IIR_out         : out signed (15 downto 0);   -- Output

	B0 : in signed(W_coef-1 downto 0);  
   B1 : in signed(W_coef-1 downto 0);
   B2 : in signed(W_coef-1 downto 0);
   A0 : in signed(W_coef-1 downto 0);
   A1 : in signed(W_coef-1 downto 0);
   A2 : in signed(W_coef-1 downto 0)
);
end component;

type cA0_array_type is array (0 to 625) of integer;  --626 length
signal A0 : cA0_array_type:=(262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144 ,262144
);

type cA1_array_type is array (0 to 625) of integer;
signal A1 : cA1_array_type:=( -509973,-509955,-509937,-509919,-509901,-509883,-509864,-509846,-509827,-509808,-509789,-509770,-509751,-509732,-509712,-509692,-509672,-509653,-509632,-509612,-509592,-509571,-509551,-509530,-509509,-509488,-509467,-509445,-509424,-509402,-509381,-509359,-509337,-509314,-509292,-509270,-509247,-509224,-509201,-509178,-509155,-509132,-509108,-509085,-509061,-509037,-509013,-508989,-508965,-508940,-508916,-508891,-508866,-508841,-508816,-508791,-508766,-508740,-508714,-508689,-508663,-508637,-508610,-508584,-508557,-508531,-508504,-508477,-508450,-508423,-508396,-508368,-508340,-508313,-508285,-508257,-508229,-508200,-508172,-508143,-508114,-508086,-508056,-508027,-507998,-507969,-507939,-507909,-507879,-507849,-507819,-507789,-507759,-507728,-507697,-507667,-507636,-507605,-507573,-507542,-507510,-507479,-507447,-507415,-507383,-507351,-507318,-507286,-507253,-507220,-507187,-507154,-507121,-507088,-507054,-507021,-506987,-506953,-506919,-506885,-506851,-506816,-506782,-506747,-506712,-506677,-506642,-506607,-506571,-506536,-506500,-506464,-506428,-506392,-506356,-506319,-506283,-506246,-506209,-506173,-506135,-506098,-506061,-506023,-505986,-505948,-505910,-505872,-505834,-505795,-505757,-505718,-505680,-505641,-505602,-505563,-505523,-505484,-505444,-505405,-505365,-505325,-505285,-505244,-505204,-505163,-505123,-505082,-505041,-505000,-504959,-504917,-504876,-504834,-504792,-504750,-504708,-504666,-504624,-504581,-504539,-504496,-504453,-504410,-504367,-504323,-504280,-504236,-504193,-504149,-504105,-504061,-504016,-503972,-503927,-503883,-503838,-503793,-503748,-503702,-503657,-503612,-503566,-503520,-503474,-503428,-503382,-503335,-503289,-503242,-503196,-503149,-503102,-503054,-503007,-502960,-502912,-502864,-502816,-502768,-502720,-502672,-502624,-502575,-502526,-502478,-502429,-502379,-502330,-502281,-502231,-502182,-502132,-502082,-502032,-501982,-501931,-501881,-501830,-501779,-501728,-501677,-501626,-501575,-501523,-501472,-501420,-501368,-501316,-501264,-501212,-501159,-501107,-501054,-501001,-500948,-500895,-500842,-500789,-500735,-500682,-500628,-500574,-500520,-500466,-500411,-500357,-500302,-500247,-500193,-500138,-500082,-500027,-499972,-499916,-499860,-499805,-499749,-499692,-499636,-499580,-499523,-499467,-499410,-499353,-499296,-499239,-499181,-499124,-499066,-499008,-498950,-498892,-498834,-498776,-498717,-498659,-498600,-498541,-498482,-498423,-498364,-498305,-498245,-498185,-498126,-498066,-498005,-497945,-497885,-497824,-497764,-497703,-497642,-497581,-497520,-497459,-497397,-497336,-497274,-497212,-497150,-497088,-497026,-496963,-496901,-496838,-496775,-496712,-496649,-496586,-496523,-496459,-496395,-496332,-496268,-496204,-496140,-496075,-496011,-495946,-495882,-495817,-495752,-495687,-495621,-495556,-495490,-495425,-495359,-495293,-495227,-495161,-495094,-495028,-494961,-494894,-494828,-494761,-494693,-494626,-494559,-494491,-494423,-494356,-494288,-494219,-494151,-494083,-494014,-493946,-493877,-493808,-493739,-493670,-493600,-493531,-493461,-493392,-493322,-493252,-493182,-493111,-493041,-492970,-492900,-492829,-492758,-492687,-492616,-492544,-492473,-492401,-492329,-492257,-492185,-492113,-492041,-491969,-491896,-491823,-491750,-491677,-491604,-491531,-491458,-491384,-491311,-491237,-491163,-491089,-491015,-490940,-490866,-490791,-490716,-490642,-490567,-490492,-490416,-490341,-490265,-490190,-490114,-490038,-489962,-489886,-489809,-489733,-489656,-489579,-489503,-489426,-489348,-489271,-489194,-489116,-489039,-488961,-488883,-488805,-488726,-488648,-488570,-488491,-488412,-488333,-488254,-488175,-488096,-488016,-487937,-487857,-487777,-487697,-487617,-487537,-487457,-487376,-487296,-487215,-487134,-487053,-486972,-486891,-486809,-486728,-486646,-486564,-486482,-486400,-486318,-486235,-486153,-486070,-485987,-485905,-485822,-485738,-485655,-485572,-485488,-485404,-485321,-485237,-485153,-485068,-484984,-484899,-484815,-484730,-484645,-484560,-484475,-484390,-484304,-484219,-484133,-484047,-483961,-483875,-483789,-483703,-483616,-483530,-483443,-483356,-483269,-483182,-483095,-483007,-482920,-482832,-482744,-482656,-482568,-482480,-482392,-482303,-482214,-482126,-482037,-481948,-481859,-481769,-481680,-481591,-481501,-481411,-481321,-481231,-481141,-481051,-480960,-480870,-480779,-480688,-480597,-480506,-480415,-480323,-480232,-480140,-480048,-479957,-479864,-479772,-479680,-479588,-479495,-479402,-479310,-479217,-479124,-479030,-478937,-478843,-478750,-478656,-478562,-478468,-478374,-478280,-478185,-478091,-477996,-477902,-477807,-477712,-477616,-477521,-477426,-477330,-477234,-477138,-477043,-476946,-476850,-476754,-476657,-476561,-476464,-476367,-476270,-476173,-476076,-475978,-475881,-475783,-475685,-475587,-475489,-475391,-475293,-475194,-475096,-474997,-474898,-474799,-474700,-474601,-474502,-474402,-474302,-474203,-474103,-474003,-473903,-473802,-473702,-473602,-473501,-473400,-473299,-473198,-473097,-472996,-472894,-472793,-472691,-472589,-472487,-472385,-472283,-472181,-472078
);

type cA2_array_type is array (0 to 625) of integer;
signal A2 : cA2_array_type:= (248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765,248765
);

type cB0_array_type is array (0 to 625) of integer;
signal B0 : cB0_array_type:= (6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689,6689
);

type cB1_array_type is array (0 to 625) of integer;
signal B1 : cB1_array_type:= (others => 0);

type cB2_array_type is array (0 to 625) of integer;
signal B2 : cB2_array_type:=(-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689,-6689
);

signal constA0 : signed(w_coef-1 downto 0):= to_signed(A0(0),w_coef);
signal constA1 : signed(w_coef-1 downto 0):= to_signed(A1(0),w_coef);
signal constA2 : signed(w_coef-1 downto 0):= to_signed(A2(0),w_coef);
signal constB0 : signed(w_coef-1 downto 0):= to_signed(B0(0),w_coef);
signal constB1 : signed(w_coef-1 downto 0):= to_signed(B1(0),w_coef);
signal constB2 : signed(w_coef-1 downto 0):= to_signed(B2(0),w_coef);

signal BP_out : signed(W_in-1 downto 0) := (others =>'0');
signal data_out_temp:  signed(W_in-1 downto 0) := (others =>'0');

begin

process(CLK_50,nReset)
variable direction: std_logic := '0';
variable counter : integer := 0;
begin
if(nReset ='0') then
	counter := 0;
elsif(rising_edge(CLK_50)) then
	if(new_val = '1') then
		data_out_temp <= BP_out+data_in; -- output 
		if(direction = '0') then
			constA0 <= to_signed(A0(counter),w_coef);
			constA1 <= to_signed(A1(counter),w_coef);
			constA2 <= to_signed(A2(counter),w_coef);
			constB0 <= to_signed(B0(counter),w_coef);
			constB1 <= to_signed(B1(counter),w_coef);
			constB2 <= to_signed(B2(counter),w_coef);
			counter := counter + 1;
			if(counter = 625) then
				direction := '1';
			end if;
		if(direction = '1') then
			constA0 <= to_signed(A0(counter),w_coef);
			constA1 <= to_signed(A1(counter),w_coef);
			constA2 <= to_signed(A2(counter),w_coef);
			constB0 <= to_signed(B0(counter),w_coef);
			constB1 <= to_signed(B1(counter),w_coef);
			constB2 <= to_signed(B2(counter),w_coef);
			counter := counter - 1;
			if (counter = 0) then
				direction := '0';
			end if;
		end if;
	end if;
end if;
end if;
end process;

IIRDF_inst : IIRDF1 
generic map(
    W_in => W_in,
	 W_coef => W_coef

)
port map(
	iCLK => CLK_50,          
	iRESET_N => nReset,      
	new_val => new_val,        
	IIR_in => data_in,                 
	IIR_out => BP_out ,        

	B0 => constB0,
   B1 => constB1,
   B2 => constB2,
   A0 => constA0,
   A1 => constA1,
   A2 => constA2
);

process(CLK_50,nReset)
begin
if nReset = '0' then
	data_out <= (others => '0');
elsif(rising_edge(CLK_50)) then
	if WahWah_EN = '0' then
		data_out <= data_in;
	elsif WahWah_EN = '1' then
		data_out <= data_out_temp + data_in;
	end if;
end if;
end process;
end;